LIBRARY ieee; 
LIBRARY std; 
USE ieee.std_logic_1164.all; 
USE ieee.std_logic_arith.all; 
USE ieee.std_logic_unsigned.all; 
USE std.textio.all; 
LIBRARY work; 
 
entity PCSystem is 
 
generic(numberOfBits : integer := 23);
port( 
v1 : in std_logic_vector (22 DOWNTO 0);
v2 : in std_logic_vector (22 DOWNTO 0);
v3 : in std_logic_vector (22 DOWNTO 0);
v4 : in std_logic_vector (22 DOWNTO 0);
v5 : in std_logic_vector (22 DOWNTO 0);
v6 : in std_logic_vector (22 DOWNTO 0);
v7 : in std_logic_vector (22 DOWNTO 0);
v8 : in std_logic_vector (22 DOWNTO 0);
v9 : in std_logic_vector (22 DOWNTO 0);
v10 : in std_logic_vector (22 DOWNTO 0);
v11 : in std_logic_vector (22 DOWNTO 0);
v12 : in std_logic_vector (22 DOWNTO 0);
v13 : in std_logic_vector (22 DOWNTO 0);
v14 : in std_logic_vector (22 DOWNTO 0);
v15 : in std_logic_vector (22 DOWNTO 0);
v16 : in std_logic_vector (22 DOWNTO 0);
vb1 : in std_logic_vector (22 DOWNTO 0);
vb2 : in std_logic_vector (22 DOWNTO 0);
vb3 : in std_logic_vector (22 DOWNTO 0);
vb4 : in std_logic_vector (22 DOWNTO 0);
vb5 : in std_logic_vector (22 DOWNTO 0);
vb6 : in std_logic_vector (22 DOWNTO 0);
vb7 : in std_logic_vector (22 DOWNTO 0);
vb8 : in std_logic_vector (22 DOWNTO 0);
vb9 : in std_logic_vector (22 DOWNTO 0);
vb10 : in std_logic_vector (22 DOWNTO 0);
vb11 : in std_logic_vector (22 DOWNTO 0);
vb12 : in std_logic_vector (22 DOWNTO 0);
vb13 : in std_logic_vector (22 DOWNTO 0);
vb14 : in std_logic_vector (22 DOWNTO 0);
vb15 : in std_logic_vector (22 DOWNTO 0);
vb16 : in std_logic_vector (22 DOWNTO 0);
vout : out std_logic_vector (22 DOWNTO 0)); 
 
end PCSystem; 

architecture rtl of PCSystem is 
 
Signal ProductNode_POSIT0weight : std_logic_vector ( 22 downto 0 ) := "00111111011111000000111";

Signal ProductNode_POSIT0Output_0: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1weight : std_logic_vector ( 22 downto 0 ) := "00111111110100011100010";

Signal ProductNode_POSIT1Output_1: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2weight : std_logic_vector ( 22 downto 0 ) := "00111111111100111010110";

Signal ProductNode_POSIT2Output_2: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3weight : std_logic_vector ( 22 downto 0 ) := "00111111101110110110111";

Signal ProductNode_POSIT3Output_3: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4weight : std_logic_vector ( 22 downto 0 ) := "00111111101111011101001";

Signal ProductNode_POSIT4Output_4: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5weight : std_logic_vector ( 22 downto 0 ) := "00111111000001000101100";

Signal ProductNode_POSIT5Output_5: std_logic_vector (22 downto 0);
Signal SumNode_POSIT0Output_6: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6Output_7: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7weight : std_logic_vector ( 22 downto 0 ) := "00111111101011111101001";

Signal ProductNode_POSIT7Output_8: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8weight : std_logic_vector ( 22 downto 0 ) := "00111111110001100000001";

Signal ProductNode_POSIT8Output_9: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9weight : std_logic_vector ( 22 downto 0 ) := "00111110111100110010000";

Signal ProductNode_POSIT9Output_10: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10weight : std_logic_vector ( 22 downto 0 ) := "00111110111001111111000";

Signal ProductNode_POSIT10Output_11: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1Output_12: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11Output_13: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT12weight : std_logic_vector ( 22 downto 0 ) := "00111111011100011010001";

Signal ProductNode_POSIT12Output_14: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT13weight : std_logic_vector ( 22 downto 0 ) := "00111111100001110010111";

Signal ProductNode_POSIT13Output_15: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2Output_16: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT14Output_17: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT15weight : std_logic_vector ( 22 downto 0 ) := "00111111001000000101101";

Signal ProductNode_POSIT15Output_18: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT16weight : std_logic_vector ( 22 downto 0 ) := "00111111110001100000001";

Signal ProductNode_POSIT16Output_19: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT17weight : std_logic_vector ( 22 downto 0 ) := "00111111110000110011011";

Signal ProductNode_POSIT17Output_20: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT18weight : std_logic_vector ( 22 downto 0 ) := "00111110111001111111000";

Signal ProductNode_POSIT18Output_21: std_logic_vector (22 downto 0);
Signal SumNode_POSIT3Output_22: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT19Output_23: std_logic_vector (22 downto 0);
Signal SumNode_POSIT4Output_24: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT20Output_25: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT21weight : std_logic_vector ( 22 downto 0 ) := "00111111000010010010001";

Signal ProductNode_POSIT21Output_26: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT25weight : std_logic_vector ( 22 downto 0 ) := "00111111010101001100011";

Signal ProductNode_POSIT25Output_31: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT26weight : std_logic_vector ( 22 downto 0 ) := "00111111010110111111101";

Signal ProductNode_POSIT26Output_32: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT27weight : std_logic_vector ( 22 downto 0 ) := "00111110001101111101000";

Signal ProductNode_POSIT27Output_33: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT28weight : std_logic_vector ( 22 downto 0 ) := "00111111100100100000001";

Signal ProductNode_POSIT28Output_34: std_logic_vector (22 downto 0);
Signal SumNode_POSIT6Output_35: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT29Output_36: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT33weight : std_logic_vector ( 22 downto 0 ) := "00111111100101011001110";

Signal ProductNode_POSIT33Output_41: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT34weight : std_logic_vector ( 22 downto 0 ) := "00111111010110111111101";

Signal ProductNode_POSIT34Output_42: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT35weight : std_logic_vector ( 22 downto 0 ) := "00111111111010010000010";

Signal ProductNode_POSIT35Output_43: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT36weight : std_logic_vector ( 22 downto 0 ) := "00111111100100100000001";

Signal ProductNode_POSIT36Output_44: std_logic_vector (22 downto 0);
Signal SumNode_POSIT8Output_45: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT37Output_46: std_logic_vector (22 downto 0);
Signal SumNode_POSIT9Output_47: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT38Output_48: std_logic_vector (22 downto 0);
Signal SumNode_POSIT10Output_49: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT39Output_50: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT40weight : std_logic_vector ( 22 downto 0 ) := "00111111110010001111101";

Signal ProductNode_POSIT40Output_51: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT41weight : std_logic_vector ( 22 downto 0 ) := "00111111101010111111011";

Signal ProductNode_POSIT41Output_52: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT42weight : std_logic_vector ( 22 downto 0 ) := "00111111100111110110110";

Signal ProductNode_POSIT42Output_53: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT43weight : std_logic_vector ( 22 downto 0 ) := "00111111101010010001010";

Signal ProductNode_POSIT43Output_54: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT44weight : std_logic_vector ( 22 downto 0 ) := "00111111111100111111010";

Signal ProductNode_POSIT44Output_55: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT45weight : std_logic_vector ( 22 downto 0 ) := "00111111001010000001001";

Signal ProductNode_POSIT45Output_56: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT46weight : std_logic_vector ( 22 downto 0 ) := "00111110001000100011001";

Signal ProductNode_POSIT46Output_57: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT47weight : std_logic_vector ( 22 downto 0 ) := "00111111001101111101010";

Signal ProductNode_POSIT47Output_58: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT48weight : std_logic_vector ( 22 downto 0 ) := "00111111110110110101110";

Signal ProductNode_POSIT48Output_59: std_logic_vector (22 downto 0);
Signal SumNode_POSIT11Output_60: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT49Output_61: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT50weight : std_logic_vector ( 22 downto 0 ) := "00111111110010110011011";

Signal ProductNode_POSIT50Output_62: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT53weight : std_logic_vector ( 22 downto 0 ) := "00111111001011011101011";

Signal ProductNode_POSIT53Output_65: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT54weight : std_logic_vector ( 22 downto 0 ) := "00111111101010110010000";

Signal ProductNode_POSIT54Output_66: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT57weight : std_logic_vector ( 22 downto 0 ) := "00111111101001000001010";

Signal ProductNode_POSIT57Output_69: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT58weight : std_logic_vector ( 22 downto 0 ) := "00111111100100010000111";

Signal ProductNode_POSIT58Output_70: std_logic_vector (22 downto 0);
Signal SumNode_POSIT12Output_71: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT59Output_72: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT60weight : std_logic_vector ( 22 downto 0 ) := "00111111001100110111010";

Signal ProductNode_POSIT60Output_73: std_logic_vector (22 downto 0);
Signal SumNode_POSIT13Output_74: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT61Output_75: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT62weight : std_logic_vector ( 22 downto 0 ) := "00111111111000110110110";

Signal ProductNode_POSIT62Output_76: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT63weight : std_logic_vector ( 22 downto 0 ) := "00111111111000111100011";

Signal ProductNode_POSIT63Output_77: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT64weight : std_logic_vector ( 22 downto 0 ) := "00111110011000011100101";

Signal ProductNode_POSIT64Output_78: std_logic_vector (22 downto 0);
Signal SumNode_POSIT14Output_79: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT65Output_80: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT66weight : std_logic_vector ( 22 downto 0 ) := "00111111111111100101100";

Signal ProductNode_POSIT66Output_81: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT67weight : std_logic_vector ( 22 downto 0 ) := "00111111000111100000001";

Signal ProductNode_POSIT67Output_82: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT68weight : std_logic_vector ( 22 downto 0 ) := "00111111101100001111111";

Signal ProductNode_POSIT68Output_83: std_logic_vector (22 downto 0);
Signal SumNode_POSIT15Output_84: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT69Output_85: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT70weight : std_logic_vector ( 22 downto 0 ) := "00111100010100111011011";

Signal ProductNode_POSIT70Output_86: std_logic_vector (22 downto 0);
Signal SumNode_POSIT16Output_87: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT71Output_88: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT72weight : std_logic_vector ( 22 downto 0 ) := "00111110110111000001011";

Signal ProductNode_POSIT72Output_89: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT73weight : std_logic_vector ( 22 downto 0 ) := "00111101111111001111110";

Signal ProductNode_POSIT73Output_90: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT74weight : std_logic_vector ( 22 downto 0 ) := "00111111101010110000011";

Signal ProductNode_POSIT74Output_91: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT75weight : std_logic_vector ( 22 downto 0 ) := "00111111110001100000011";

Signal ProductNode_POSIT75Output_92: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT76weight : std_logic_vector ( 22 downto 0 ) := "00111111111101110000011";

Signal ProductNode_POSIT76Output_93: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT77weight : std_logic_vector ( 22 downto 0 ) := "00111111111100000011000";

Signal ProductNode_POSIT77Output_94: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT78weight : std_logic_vector ( 22 downto 0 ) := "00111101000110010111001";

Signal ProductNode_POSIT78Output_95: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT79weight : std_logic_vector ( 22 downto 0 ) := "00111111000110101000001";

Signal ProductNode_POSIT79Output_96: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT80weight : std_logic_vector ( 22 downto 0 ) := "00111111101111001000100";

Signal ProductNode_POSIT80Output_97: std_logic_vector (22 downto 0);
Signal SumNode_POSIT17Output_98: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT81Output_99: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT82weight : std_logic_vector ( 22 downto 0 ) := "00111111110010110011011";

Signal ProductNode_POSIT82Output_100: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT85weight : std_logic_vector ( 22 downto 0 ) := "00111110111001111110011";

Signal ProductNode_POSIT85Output_103: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT86weight : std_logic_vector ( 22 downto 0 ) := "00111111101011111011011";

Signal ProductNode_POSIT86Output_104: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT89weight : std_logic_vector ( 22 downto 0 ) := "00111111101100101011111";

Signal ProductNode_POSIT89Output_107: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT90weight : std_logic_vector ( 22 downto 0 ) := "00111111100000000000000";

Signal ProductNode_POSIT90Output_108: std_logic_vector (22 downto 0);
Signal SumNode_POSIT18Output_109: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT91Output_110: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT92weight : std_logic_vector ( 22 downto 0 ) := "00111111001100110111010";

Signal ProductNode_POSIT92Output_111: std_logic_vector (22 downto 0);
Signal SumNode_POSIT19Output_112: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT93Output_113: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT94weight : std_logic_vector ( 22 downto 0 ) := "00111111101100111001011";

Signal ProductNode_POSIT94Output_114: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT98weight : std_logic_vector ( 22 downto 0 ) := "00111111111110010011111";

Signal ProductNode_POSIT98Output_119: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT102weight : std_logic_vector ( 22 downto 0 ) := "00111101010110000001110";

Signal ProductNode_POSIT102Output_124: std_logic_vector (22 downto 0);
Signal SumNode_POSIT22Output_125: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT103Output_126: std_logic_vector (22 downto 0);
Signal SumNode_POSIT23Output_127: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT104Output_128: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT105weight : std_logic_vector ( 22 downto 0 ) := "00111110101100011000011";

Signal ProductNode_POSIT105Output_129: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT106weight : std_logic_vector ( 22 downto 0 ) := "00111111101111111110110";

Signal ProductNode_POSIT106Output_130: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT112weight : std_logic_vector ( 22 downto 0 ) := "00111111100101011011010";

Signal ProductNode_POSIT112Output_137: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT114weight : std_logic_vector ( 22 downto 0 ) := "00111111010101001001010";

Signal ProductNode_POSIT114Output_139: std_logic_vector (22 downto 0);
Signal SumNode_POSIT25Output_140: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT115Output_141: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT120weight : std_logic_vector ( 22 downto 0 ) := "00111111100101011011010";

Signal ProductNode_POSIT120Output_147: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT122weight : std_logic_vector ( 22 downto 0 ) := "00111111010101001001010";

Signal ProductNode_POSIT122Output_149: std_logic_vector (22 downto 0);
Signal SumNode_POSIT27Output_150: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT123Output_151: std_logic_vector (22 downto 0);
Signal SumNode_POSIT28Output_152: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT124Output_153: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT130weight : std_logic_vector ( 22 downto 0 ) := "00111111000010010111010";

Signal ProductNode_POSIT130Output_160: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT132weight : std_logic_vector ( 22 downto 0 ) := "00111111101110110100010";

Signal ProductNode_POSIT132Output_162: std_logic_vector (22 downto 0);
Signal SumNode_POSIT30Output_163: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT133Output_164: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT138weight : std_logic_vector ( 22 downto 0 ) := "00111111000010010111010";

Signal ProductNode_POSIT138Output_170: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT140weight : std_logic_vector ( 22 downto 0 ) := "00111111101110110100010";

Signal ProductNode_POSIT140Output_172: std_logic_vector (22 downto 0);
Signal SumNode_POSIT32Output_173: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT141Output_174: std_logic_vector (22 downto 0);
Signal SumNode_POSIT33Output_175: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT142Output_176: std_logic_vector (22 downto 0);
Signal SumNode_POSIT34Output_177: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT143Output_178: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT166weight : std_logic_vector ( 22 downto 0 ) := "00111110011001001001101";

Signal ProductNode_POSIT166Output_204: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT170weight : std_logic_vector ( 22 downto 0 ) := "00111111111111100101101";

Signal ProductNode_POSIT170Output_209: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT174weight : std_logic_vector ( 22 downto 0 ) := "00111100010100101001100";

Signal ProductNode_POSIT174Output_214: std_logic_vector (22 downto 0);
Signal SumNode_POSIT40Output_215: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT175Output_216: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT198weight : std_logic_vector ( 22 downto 0 ) := "00111111000110001101000";

Signal ProductNode_POSIT198Output_242: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT202weight : std_logic_vector ( 22 downto 0 ) := "00111111111111111101111";

Signal ProductNode_POSIT202Output_247: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT206weight : std_logic_vector ( 22 downto 0 ) := "00111010100001000001111";

Signal ProductNode_POSIT206Output_252: std_logic_vector (22 downto 0);
Signal SumNode_POSIT46Output_253: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT207Output_254: std_logic_vector (22 downto 0);
Signal SumNode_POSIT47Output_255: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT208Output_256: std_logic_vector (22 downto 0);
Signal SumNode_POSIT48Output_257: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT209Output_258: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT211weight : std_logic_vector ( 22 downto 0 ) := "00111101110001010010100";

Signal ProductNode_POSIT211Output_260: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT248Output_308: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT272weight : std_logic_vector ( 22 downto 0 ) := "00111111001101110011110";

Signal ProductNode_POSIT272Output_335: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT273weight : std_logic_vector ( 22 downto 0 ) := "00111111101001000110000";

Signal ProductNode_POSIT273Output_336: std_logic_vector (22 downto 0);
Signal SumNode_POSIT63Output_337: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT274Output_338: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT275weight : std_logic_vector ( 22 downto 0 ) := "00111111111001011010011";

Signal ProductNode_POSIT275Output_339: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT276weight : std_logic_vector ( 22 downto 0 ) := "00111011111000011111011";

Signal ProductNode_POSIT276Output_340: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT277weight : std_logic_vector ( 22 downto 0 ) := "00111111111111110001111";

Signal ProductNode_POSIT277Output_341: std_logic_vector (22 downto 0);
Signal SumNode_POSIT64Output_342: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT278Output_343: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT279weight : std_logic_vector ( 22 downto 0 ) := "00111110010100101100100";

Signal ProductNode_POSIT279Output_344: std_logic_vector (22 downto 0);
Signal SumNode_POSIT65Output_345: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT280Output_346: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT307weight : std_logic_vector ( 22 downto 0 ) := "00111111110100111101100";

Signal ProductNode_POSIT307Output_377: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT311weight : std_logic_vector ( 22 downto 0 ) := "00111110101100001001110";

Signal ProductNode_POSIT311Output_382: std_logic_vector (22 downto 0);
Signal SumNode_POSIT71Output_383: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT312Output_384: std_logic_vector (22 downto 0);
Signal SumNode_POSIT72Output_385: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT313Output_386: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT315weight : std_logic_vector ( 22 downto 0 ) := "00111111000000000010010";

Signal ProductNode_POSIT315Output_388: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT352Output_436: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT379weight : std_logic_vector ( 22 downto 0 ) := "00111111110010101000000";

Signal ProductNode_POSIT379Output_467: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT383weight : std_logic_vector ( 22 downto 0 ) := "00111110110101011111111";

Signal ProductNode_POSIT383Output_472: std_logic_vector (22 downto 0);
Signal SumNode_POSIT89Output_473: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT384Output_474: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT411weight : std_logic_vector ( 22 downto 0 ) := "00111111101101101101100";

Signal ProductNode_POSIT411Output_505: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT415weight : std_logic_vector ( 22 downto 0 ) := "00111111000100100100111";

Signal ProductNode_POSIT415Output_510: std_logic_vector (22 downto 0);
Signal SumNode_POSIT95Output_511: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT416Output_512: std_logic_vector (22 downto 0);
Signal SumNode_POSIT96Output_513: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT417Output_514: std_logic_vector (22 downto 0);
Signal SumNode_POSIT97Output_515: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT418Output_516: std_logic_vector (22 downto 0);
Signal SumNode_POSIT98Output_517: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT419Output_518: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT422weight : std_logic_vector ( 22 downto 0 ) := "00111111011111001111111";

Signal ProductNode_POSIT422Output_521: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT439Output_543: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT440weight : std_logic_vector ( 22 downto 0 ) := "00111111100000011000000";

Signal ProductNode_POSIT440Output_544: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT457Output_566: std_logic_vector (22 downto 0);
Signal SumNode_POSIT109Output_567: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT458Output_568: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT463weight : std_logic_vector ( 22 downto 0 ) := "00111101110000001010100";

Signal ProductNode_POSIT463Output_573: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT467weight : std_logic_vector ( 22 downto 0 ) := "00111110100100101000111";

Signal ProductNode_POSIT467Output_577: std_logic_vector (22 downto 0);
Signal SumNode_POSIT110Output_578: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT468Output_579: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT469weight : std_logic_vector ( 22 downto 0 ) := "00111110111011010001001";

Signal ProductNode_POSIT469Output_580: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT473weight : std_logic_vector ( 22 downto 0 ) := "00111111001010011011110";

Signal ProductNode_POSIT473Output_584: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT477weight : std_logic_vector ( 22 downto 0 ) := "00111111010111011110000";

Signal ProductNode_POSIT477Output_588: std_logic_vector (22 downto 0);
Signal SumNode_POSIT111Output_589: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT478Output_590: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT479weight : std_logic_vector ( 22 downto 0 ) := "00111110001110010000011";

Signal ProductNode_POSIT479Output_591: std_logic_vector (22 downto 0);
Signal SumNode_POSIT112Output_592: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT480Output_593: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT481weight : std_logic_vector ( 22 downto 0 ) := "00111111101111011010100";

Signal ProductNode_POSIT481Output_594: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT485weight : std_logic_vector ( 22 downto 0 ) := "00111111111110000111011";

Signal ProductNode_POSIT485Output_599: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT489weight : std_logic_vector ( 22 downto 0 ) := "00111101011100010001110";

Signal ProductNode_POSIT489Output_604: std_logic_vector (22 downto 0);
Signal SumNode_POSIT115Output_605: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT490Output_606: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT495weight : std_logic_vector ( 22 downto 0 ) := "00111101100011111001110";

Signal ProductNode_POSIT495Output_611: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT499weight : std_logic_vector ( 22 downto 0 ) := "00111111000001101110111";

Signal ProductNode_POSIT499Output_615: std_logic_vector (22 downto 0);
Signal SumNode_POSIT116Output_616: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT500Output_617: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT501weight : std_logic_vector ( 22 downto 0 ) := "00111110111011010001001";

Signal ProductNode_POSIT501Output_618: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT505weight : std_logic_vector ( 22 downto 0 ) := "00111111001000001001000";

Signal ProductNode_POSIT505Output_622: std_logic_vector (22 downto 0);
Signal SumNode_POSIT117Output_627: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT510Output_628: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT511weight : std_logic_vector ( 22 downto 0 ) := "00111110001110010000011";

Signal ProductNode_POSIT511Output_629: std_logic_vector (22 downto 0);
Signal SumNode_POSIT118Output_630: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT512Output_631: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT513weight : std_logic_vector ( 22 downto 0 ) := "00111111100101000101011";

Signal ProductNode_POSIT513Output_632: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT517weight : std_logic_vector ( 22 downto 0 ) := "00111111111010100100111";

Signal ProductNode_POSIT517Output_637: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT521weight : std_logic_vector ( 22 downto 0 ) := "00111110001011011000011";

Signal ProductNode_POSIT521Output_642: std_logic_vector (22 downto 0);
Signal SumNode_POSIT121Output_643: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT522Output_644: std_logic_vector (22 downto 0);
Signal SumNode_POSIT122Output_645: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT523Output_646: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT543Output_671: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT561Output_694: std_logic_vector (22 downto 0);
Signal SumNode_POSIT133Output_695: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT562Output_696: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT585weight : std_logic_vector ( 22 downto 0 ) := "00111111000001001010110";

Signal ProductNode_POSIT585Output_722: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT589weight : std_logic_vector ( 22 downto 0 ) := "00111111110101101110000";

Signal ProductNode_POSIT589Output_727: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT593weight : std_logic_vector ( 22 downto 0 ) := "00111110101001000111101";

Signal ProductNode_POSIT593Output_732: std_logic_vector (22 downto 0);
Signal SumNode_POSIT139Output_733: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT594Output_734: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT617weight : std_logic_vector ( 22 downto 0 ) := "00111111010101110101001";

Signal ProductNode_POSIT617Output_760: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT621weight : std_logic_vector ( 22 downto 0 ) := "00111111111000011101001";

Signal ProductNode_POSIT621Output_765: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT625weight : std_logic_vector ( 22 downto 0 ) := "00111110011100010110101";

Signal ProductNode_POSIT625Output_770: std_logic_vector (22 downto 0);
Signal SumNode_POSIT145Output_771: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT626Output_772: std_logic_vector (22 downto 0);
Signal SumNode_POSIT146Output_773: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT627Output_774: std_logic_vector (22 downto 0);
Signal SumNode_POSIT147Output_775: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT628Output_776: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT667Output_826: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT694weight : std_logic_vector ( 22 downto 0 ) := "00111111110010101111110";

Signal ProductNode_POSIT694Output_857: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT698weight : std_logic_vector ( 22 downto 0 ) := "00111110110101000000100";

Signal ProductNode_POSIT698Output_862: std_logic_vector (22 downto 0);
Signal SumNode_POSIT164Output_863: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT699Output_864: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT726weight : std_logic_vector ( 22 downto 0 ) := "00111111101100011011010";

Signal ProductNode_POSIT726Output_895: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT730weight : std_logic_vector ( 22 downto 0 ) := "00111111000111001001011";

Signal ProductNode_POSIT730Output_900: std_logic_vector (22 downto 0);
Signal SumNode_POSIT170Output_901: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT731Output_902: std_logic_vector (22 downto 0);
Signal SumNode_POSIT171Output_903: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT732Output_904: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT771Output_954: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT798weight : std_logic_vector ( 22 downto 0 ) := "00111111101100100011100";

Signal ProductNode_POSIT798Output_985: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT802weight : std_logic_vector ( 22 downto 0 ) := "00111111000110111000110";

Signal ProductNode_POSIT802Output_990: std_logic_vector (22 downto 0);
Signal SumNode_POSIT188Output_991: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT803Output_992: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT830weight : std_logic_vector ( 22 downto 0 ) := "00111111100001101001010";

Signal ProductNode_POSIT830Output_1023: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT834weight : std_logic_vector ( 22 downto 0 ) := "00111111011100101101011";

Signal ProductNode_POSIT834Output_1028: std_logic_vector (22 downto 0);
Signal SumNode_POSIT194Output_1029: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT835Output_1030: std_logic_vector (22 downto 0);
Signal SumNode_POSIT195Output_1031: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT836Output_1032: std_logic_vector (22 downto 0);
Signal SumNode_POSIT196Output_1033: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT837Output_1034: std_logic_vector (22 downto 0);
Signal SumNode_POSIT197Output_1035: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT838Output_1036: std_logic_vector (22 downto 0);
Signal SumNode_POSIT198Output_1037: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT839Output_1038: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT840weight : std_logic_vector ( 22 downto 0 ) := "00111111001000011101010";

Signal ProductNode_POSIT840Output_1039: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT841weight : std_logic_vector ( 22 downto 0 ) := "00111111111100111010110";

Signal ProductNode_POSIT841Output_1040: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT842weight : std_logic_vector ( 22 downto 0 ) := "00111111010101011110100";

Signal ProductNode_POSIT842Output_1041: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT843weight : std_logic_vector ( 22 downto 0 ) := "00111110101010101101001";

Signal ProductNode_POSIT843Output_1042: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT844weight : std_logic_vector ( 22 downto 0 ) := "00111111110101010100101";

Signal ProductNode_POSIT844Output_1043: std_logic_vector (22 downto 0);
Signal SumNode_POSIT199Output_1044: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT845Output_1045: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT850Output_1051: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT851weight : std_logic_vector ( 22 downto 0 ) := "00111110001010011111000";

Signal ProductNode_POSIT851Output_1052: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT852weight : std_logic_vector ( 22 downto 0 ) := "00111111111010101100000";

Signal ProductNode_POSIT852Output_1053: std_logic_vector (22 downto 0);
Signal SumNode_POSIT201Output_1054: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT853Output_1055: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT858Output_1061: std_logic_vector (22 downto 0);
Signal SumNode_POSIT203Output_1062: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT859Output_1063: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT860weight : std_logic_vector ( 22 downto 0 ) := "00111111100101010000101";

Signal ProductNode_POSIT860Output_1064: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT868Output_1074: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT876Output_1084: std_logic_vector (22 downto 0);
Signal SumNode_POSIT208Output_1085: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT877Output_1086: std_logic_vector (22 downto 0);
Signal SumNode_POSIT209Output_1087: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT878Output_1088: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT889weight : std_logic_vector ( 22 downto 0 ) := "00111110110100110010000";

Signal ProductNode_POSIT889Output_1100: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT899weight : std_logic_vector ( 22 downto 0 ) := "00111111101001100100010";

Signal ProductNode_POSIT899Output_1111: std_logic_vector (22 downto 0);
Signal SumNode_POSIT212Output_1112: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT900Output_1113: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT901weight : std_logic_vector ( 22 downto 0 ) := "00111111111000110110110";

Signal ProductNode_POSIT901Output_1114: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT902weight : std_logic_vector ( 22 downto 0 ) := "00111111100111000100100";

Signal ProductNode_POSIT902Output_1115: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT903weight : std_logic_vector ( 22 downto 0 ) := "00111111010001110110110";

Signal ProductNode_POSIT903Output_1116: std_logic_vector (22 downto 0);
Signal SumNode_POSIT213Output_1117: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT904Output_1118: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT905weight : std_logic_vector ( 22 downto 0 ) := "00111111111111100101100";

Signal ProductNode_POSIT905Output_1119: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT906weight : std_logic_vector ( 22 downto 0 ) := "00111110000010100110000";

Signal ProductNode_POSIT906Output_1120: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT907weight : std_logic_vector ( 22 downto 0 ) := "00111111111011101011001";

Signal ProductNode_POSIT907Output_1121: std_logic_vector (22 downto 0);
Signal SumNode_POSIT214Output_1122: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT908Output_1123: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT909weight : std_logic_vector ( 22 downto 0 ) := "00111100010100111011011";

Signal ProductNode_POSIT909Output_1124: std_logic_vector (22 downto 0);
Signal SumNode_POSIT215Output_1125: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT910Output_1126: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT921weight : std_logic_vector ( 22 downto 0 ) := "00111110110100110010000";

Signal ProductNode_POSIT921Output_1138: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT931weight : std_logic_vector ( 22 downto 0 ) := "00111111101001100100010";

Signal ProductNode_POSIT931Output_1149: std_logic_vector (22 downto 0);
Signal SumNode_POSIT218Output_1150: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT932Output_1151: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT933weight : std_logic_vector ( 22 downto 0 ) := "00111111101100111001011";

Signal ProductNode_POSIT933Output_1152: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT937weight : std_logic_vector ( 22 downto 0 ) := "00111111111110010011111";

Signal ProductNode_POSIT937Output_1157: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT941weight : std_logic_vector ( 22 downto 0 ) := "00111101010110000001110";

Signal ProductNode_POSIT941Output_1162: std_logic_vector (22 downto 0);
Signal SumNode_POSIT221Output_1163: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT942Output_1164: std_logic_vector (22 downto 0);
Signal SumNode_POSIT222Output_1165: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT943Output_1166: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT944weight : std_logic_vector ( 22 downto 0 ) := "00111101001110110100001";

Signal ProductNode_POSIT944Output_1167: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT945weight : std_logic_vector ( 22 downto 0 ) := "00111111101111111110110";

Signal ProductNode_POSIT945Output_1168: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT954Output_1179: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT962Output_1189: std_logic_vector (22 downto 0);
Signal SumNode_POSIT227Output_1190: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT963Output_1191: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT972Output_1202: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT980Output_1212: std_logic_vector (22 downto 0);
Signal SumNode_POSIT232Output_1213: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT981Output_1214: std_logic_vector (22 downto 0);
Signal SumNode_POSIT233Output_1215: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT982Output_1216: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1005weight : std_logic_vector ( 22 downto 0 ) := "00111110011001001001101";

Signal ProductNode_POSIT1005Output_1242: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1009weight : std_logic_vector ( 22 downto 0 ) := "00111111111111100101101";

Signal ProductNode_POSIT1009Output_1247: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1013weight : std_logic_vector ( 22 downto 0 ) := "00111100010100101001100";

Signal ProductNode_POSIT1013Output_1252: std_logic_vector (22 downto 0);
Signal SumNode_POSIT239Output_1253: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1014Output_1254: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1037weight : std_logic_vector ( 22 downto 0 ) := "00111111000110001101000";

Signal ProductNode_POSIT1037Output_1280: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1041weight : std_logic_vector ( 22 downto 0 ) := "00111111111111111101111";

Signal ProductNode_POSIT1041Output_1285: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1045weight : std_logic_vector ( 22 downto 0 ) := "00111010100001000001111";

Signal ProductNode_POSIT1045Output_1290: std_logic_vector (22 downto 0);
Signal SumNode_POSIT245Output_1291: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1046Output_1292: std_logic_vector (22 downto 0);
Signal SumNode_POSIT246Output_1293: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1047Output_1294: std_logic_vector (22 downto 0);
Signal SumNode_POSIT247Output_1295: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1048Output_1296: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1050weight : std_logic_vector ( 22 downto 0 ) := "00111101110001010010100";

Signal ProductNode_POSIT1050Output_1298: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1087Output_1346: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1111weight : std_logic_vector ( 22 downto 0 ) := "00111110100110001101101";

Signal ProductNode_POSIT1111Output_1373: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1112weight : std_logic_vector ( 22 downto 0 ) := "00111111110110011100100";

Signal ProductNode_POSIT1112Output_1374: std_logic_vector (22 downto 0);
Signal SumNode_POSIT262Output_1375: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1113Output_1376: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1114weight : std_logic_vector ( 22 downto 0 ) := "00111111111001011010011";

Signal ProductNode_POSIT1114Output_1377: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1115weight : std_logic_vector ( 22 downto 0 ) := "00111010101110011101110";

Signal ProductNode_POSIT1115Output_1378: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1116weight : std_logic_vector ( 22 downto 0 ) := "00111111111111111101000";

Signal ProductNode_POSIT1116Output_1379: std_logic_vector (22 downto 0);
Signal SumNode_POSIT263Output_1380: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1117Output_1381: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1118weight : std_logic_vector ( 22 downto 0 ) := "00111110010100101100100";

Signal ProductNode_POSIT1118Output_1382: std_logic_vector (22 downto 0);
Signal SumNode_POSIT264Output_1383: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1119Output_1384: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1146weight : std_logic_vector ( 22 downto 0 ) := "00111111110100111101100";

Signal ProductNode_POSIT1146Output_1415: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1150weight : std_logic_vector ( 22 downto 0 ) := "00111110101100001001110";

Signal ProductNode_POSIT1150Output_1420: std_logic_vector (22 downto 0);
Signal SumNode_POSIT270Output_1421: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1151Output_1422: std_logic_vector (22 downto 0);
Signal SumNode_POSIT271Output_1423: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1152Output_1424: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1154weight : std_logic_vector ( 22 downto 0 ) := "00111111000000000010010";

Signal ProductNode_POSIT1154Output_1426: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1191Output_1474: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1218weight : std_logic_vector ( 22 downto 0 ) := "00111111110010101000000";

Signal ProductNode_POSIT1218Output_1505: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1222weight : std_logic_vector ( 22 downto 0 ) := "00111110110101011111111";

Signal ProductNode_POSIT1222Output_1510: std_logic_vector (22 downto 0);
Signal SumNode_POSIT288Output_1511: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1223Output_1512: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1250weight : std_logic_vector ( 22 downto 0 ) := "00111111101101101101100";

Signal ProductNode_POSIT1250Output_1543: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1254weight : std_logic_vector ( 22 downto 0 ) := "00111111000100100100111";

Signal ProductNode_POSIT1254Output_1548: std_logic_vector (22 downto 0);
Signal SumNode_POSIT294Output_1549: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1255Output_1550: std_logic_vector (22 downto 0);
Signal SumNode_POSIT295Output_1551: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1256Output_1552: std_logic_vector (22 downto 0);
Signal SumNode_POSIT296Output_1553: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1257Output_1554: std_logic_vector (22 downto 0);
Signal SumNode_POSIT297Output_1555: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1258Output_1556: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1261weight : std_logic_vector ( 22 downto 0 ) := "00111111001101010110111";

Signal ProductNode_POSIT1261Output_1559: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1278Output_1581: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1279weight : std_logic_vector ( 22 downto 0 ) := "00111111101001010100100";

Signal ProductNode_POSIT1279Output_1582: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1296Output_1604: std_logic_vector (22 downto 0);
Signal SumNode_POSIT308Output_1605: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1297Output_1606: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1308weight : std_logic_vector ( 22 downto 0 ) := "00111111110001001011101";

Signal ProductNode_POSIT1308Output_1618: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1318weight : std_logic_vector ( 22 downto 0 ) := "00111111111010001101111";

Signal ProductNode_POSIT1318Output_1629: std_logic_vector (22 downto 0);
Signal SumNode_POSIT311Output_1630: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1319Output_1631: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1320weight : std_logic_vector ( 22 downto 0 ) := "00111111101111011010100";

Signal ProductNode_POSIT1320Output_1632: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1324weight : std_logic_vector ( 22 downto 0 ) := "00111111111110000111011";

Signal ProductNode_POSIT1324Output_1637: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1328weight : std_logic_vector ( 22 downto 0 ) := "00111101011100010001110";

Signal ProductNode_POSIT1328Output_1642: std_logic_vector (22 downto 0);
Signal SumNode_POSIT314Output_1643: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1329Output_1644: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1340weight : std_logic_vector ( 22 downto 0 ) := "00111111110001001011101";

Signal ProductNode_POSIT1340Output_1656: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1350weight : std_logic_vector ( 22 downto 0 ) := "00111111111010001101111";

Signal ProductNode_POSIT1350Output_1667: std_logic_vector (22 downto 0);
Signal SumNode_POSIT317Output_1668: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1351Output_1669: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1352weight : std_logic_vector ( 22 downto 0 ) := "00111111100101000101011";

Signal ProductNode_POSIT1352Output_1670: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1356weight : std_logic_vector ( 22 downto 0 ) := "00111111111010100100111";

Signal ProductNode_POSIT1356Output_1675: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1360weight : std_logic_vector ( 22 downto 0 ) := "00111110001011011000011";

Signal ProductNode_POSIT1360Output_1680: std_logic_vector (22 downto 0);
Signal SumNode_POSIT320Output_1681: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1361Output_1682: std_logic_vector (22 downto 0);
Signal SumNode_POSIT321Output_1683: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1362Output_1684: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1382Output_1709: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1400Output_1732: std_logic_vector (22 downto 0);
Signal SumNode_POSIT332Output_1733: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1401Output_1734: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1424weight : std_logic_vector ( 22 downto 0 ) := "00111111000001001010110";

Signal ProductNode_POSIT1424Output_1760: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1428weight : std_logic_vector ( 22 downto 0 ) := "00111111110101101110000";

Signal ProductNode_POSIT1428Output_1765: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1432weight : std_logic_vector ( 22 downto 0 ) := "00111110101001000111101";

Signal ProductNode_POSIT1432Output_1770: std_logic_vector (22 downto 0);
Signal SumNode_POSIT338Output_1771: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1433Output_1772: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1456weight : std_logic_vector ( 22 downto 0 ) := "00111111010101110101001";

Signal ProductNode_POSIT1456Output_1798: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1460weight : std_logic_vector ( 22 downto 0 ) := "00111111111000011101001";

Signal ProductNode_POSIT1460Output_1803: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1464weight : std_logic_vector ( 22 downto 0 ) := "00111110011100010110101";

Signal ProductNode_POSIT1464Output_1808: std_logic_vector (22 downto 0);
Signal SumNode_POSIT344Output_1809: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1465Output_1810: std_logic_vector (22 downto 0);
Signal SumNode_POSIT345Output_1811: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1466Output_1812: std_logic_vector (22 downto 0);
Signal SumNode_POSIT346Output_1813: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1467Output_1814: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1506Output_1864: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1533weight : std_logic_vector ( 22 downto 0 ) := "00111111110010101111110";

Signal ProductNode_POSIT1533Output_1895: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1537weight : std_logic_vector ( 22 downto 0 ) := "00111110110101000000100";

Signal ProductNode_POSIT1537Output_1900: std_logic_vector (22 downto 0);
Signal SumNode_POSIT363Output_1901: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1538Output_1902: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1565weight : std_logic_vector ( 22 downto 0 ) := "00111111101100011011010";

Signal ProductNode_POSIT1565Output_1933: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1569weight : std_logic_vector ( 22 downto 0 ) := "00111111000111001001011";

Signal ProductNode_POSIT1569Output_1938: std_logic_vector (22 downto 0);
Signal SumNode_POSIT369Output_1939: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1570Output_1940: std_logic_vector (22 downto 0);
Signal SumNode_POSIT370Output_1941: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1571Output_1942: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1610Output_1992: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1637weight : std_logic_vector ( 22 downto 0 ) := "00111111101100100011100";

Signal ProductNode_POSIT1637Output_2023: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1641weight : std_logic_vector ( 22 downto 0 ) := "00111111000110111000110";

Signal ProductNode_POSIT1641Output_2028: std_logic_vector (22 downto 0);
Signal SumNode_POSIT387Output_2029: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1642Output_2030: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1669weight : std_logic_vector ( 22 downto 0 ) := "00111111100001101001010";

Signal ProductNode_POSIT1669Output_2061: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1673weight : std_logic_vector ( 22 downto 0 ) := "00111111011100101101011";

Signal ProductNode_POSIT1673Output_2066: std_logic_vector (22 downto 0);
Signal SumNode_POSIT393Output_2067: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1674Output_2068: std_logic_vector (22 downto 0);
Signal SumNode_POSIT394Output_2069: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1675Output_2070: std_logic_vector (22 downto 0);
Signal SumNode_POSIT395Output_2071: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1676Output_2072: std_logic_vector (22 downto 0);
Signal SumNode_POSIT396Output_2073: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1677Output_2074: std_logic_vector (22 downto 0);
Signal SumNode_POSIT397Output_2075: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1678Output_2076: std_logic_vector (22 downto 0);
Signal SumNode_POSIT398Output_2077: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1679Output_2078: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1680weight : std_logic_vector ( 22 downto 0 ) := "00111110101110001110100";

Signal ProductNode_POSIT1680Output_2079: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1681weight : std_logic_vector ( 22 downto 0 ) := "00111111100010010001111";

Signal ProductNode_POSIT1681Output_2080: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1682weight : std_logic_vector ( 22 downto 0 ) := "00111111000100000111011";

Signal ProductNode_POSIT1682Output_2081: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1683weight : std_logic_vector ( 22 downto 0 ) := "00111111010101010110000";

Signal ProductNode_POSIT1683Output_2082: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1684weight : std_logic_vector ( 22 downto 0 ) := "00111111100101010100111";

Signal ProductNode_POSIT1684Output_2083: std_logic_vector (22 downto 0);
Signal SumNode_POSIT399Output_2084: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1685Output_2085: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1686weight : std_logic_vector ( 22 downto 0 ) := "00111111001011111011001";

Signal ProductNode_POSIT1686Output_2086: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1687weight : std_logic_vector ( 22 downto 0 ) := "00111111011110010011110";

Signal ProductNode_POSIT1687Output_2087: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1688weight : std_logic_vector ( 22 downto 0 ) := "00111110010000001100001";

Signal ProductNode_POSIT1688Output_2088: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1689weight : std_logic_vector ( 22 downto 0 ) := "00111111100000110110000";

Signal ProductNode_POSIT1689Output_2089: std_logic_vector (22 downto 0);
Signal SumNode_POSIT400Output_2090: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1690Output_2091: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1691weight : std_logic_vector ( 22 downto 0 ) := "00111111000111101110100";

Signal ProductNode_POSIT1691Output_2092: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1692weight : std_logic_vector ( 22 downto 0 ) := "00111111101100001000101";

Signal ProductNode_POSIT1692Output_2093: std_logic_vector (22 downto 0);
Signal SumNode_POSIT401Output_2094: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1693Output_2095: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1694weight : std_logic_vector ( 22 downto 0 ) := "00111111101010000010011";

Signal ProductNode_POSIT1694Output_2096: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1695weight : std_logic_vector ( 22 downto 0 ) := "00111111011110010011110";

Signal ProductNode_POSIT1695Output_2097: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1696weight : std_logic_vector ( 22 downto 0 ) := "00111111111001111110011";

Signal ProductNode_POSIT1696Output_2098: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1697weight : std_logic_vector ( 22 downto 0 ) := "00111111100000110110000";

Signal ProductNode_POSIT1697Output_2099: std_logic_vector (22 downto 0);
Signal SumNode_POSIT402Output_2100: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1698Output_2101: std_logic_vector (22 downto 0);
Signal SumNode_POSIT403Output_2102: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1699Output_2103: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1700weight : std_logic_vector ( 22 downto 0 ) := "00111111101101111100010";

Signal ProductNode_POSIT1700Output_2104: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1704weight : std_logic_vector ( 22 downto 0 ) := "00111110100101111111100";

Signal ProductNode_POSIT1704Output_2109: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1705weight : std_logic_vector ( 22 downto 0 ) := "00111110110100110111100";

Signal ProductNode_POSIT1705Output_2110: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1706weight : std_logic_vector ( 22 downto 0 ) := "00111101010101110001100";

Signal ProductNode_POSIT1706Output_2111: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1707weight : std_logic_vector ( 22 downto 0 ) := "00111111110010110010000";

Signal ProductNode_POSIT1707Output_2112: std_logic_vector (22 downto 0);
Signal SumNode_POSIT405Output_2113: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1708Output_2114: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1712weight : std_logic_vector ( 22 downto 0 ) := "00111111110110100000000";

Signal ProductNode_POSIT1712Output_2119: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1713weight : std_logic_vector ( 22 downto 0 ) := "00111110110100110111100";

Signal ProductNode_POSIT1713Output_2120: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1714weight : std_logic_vector ( 22 downto 0 ) := "00111111111110010100011";

Signal ProductNode_POSIT1714Output_2121: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1715weight : std_logic_vector ( 22 downto 0 ) := "00111111110010110010000";

Signal ProductNode_POSIT1715Output_2122: std_logic_vector (22 downto 0);
Signal SumNode_POSIT407Output_2123: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1716Output_2124: std_logic_vector (22 downto 0);
Signal SumNode_POSIT408Output_2125: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1717Output_2126: std_logic_vector (22 downto 0);
Signal SumNode_POSIT409Output_2127: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1718Output_2128: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1742weight : std_logic_vector ( 22 downto 0 ) := "00111111010000110000111";

Signal ProductNode_POSIT1742Output_2155: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1743weight : std_logic_vector ( 22 downto 0 ) := "00111111100111100111100";

Signal ProductNode_POSIT1743Output_2156: std_logic_vector (22 downto 0);
Signal SumNode_POSIT413Output_2157: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1744Output_2158: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1745weight : std_logic_vector ( 22 downto 0 ) := "00111111111111100101100";

Signal ProductNode_POSIT1745Output_2159: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1749weight : std_logic_vector ( 22 downto 0 ) := "00111100010100111011011";

Signal ProductNode_POSIT1749Output_2164: std_logic_vector (22 downto 0);
Signal SumNode_POSIT415Output_2165: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1750Output_2166: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1777weight : std_logic_vector ( 22 downto 0 ) := "00111111111110010011111";

Signal ProductNode_POSIT1777Output_2197: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1781weight : std_logic_vector ( 22 downto 0 ) := "00111101010110000001110";

Signal ProductNode_POSIT1781Output_2202: std_logic_vector (22 downto 0);
Signal SumNode_POSIT421Output_2203: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1782Output_2204: std_logic_vector (22 downto 0);
Signal SumNode_POSIT422Output_2205: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1783Output_2206: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1784weight : std_logic_vector ( 22 downto 0 ) := "00111111110100111001111";

Signal ProductNode_POSIT1784Output_2207: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1785weight : std_logic_vector ( 22 downto 0 ) := "00111111000100001101101";

Signal ProductNode_POSIT1785Output_2208: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1791weight : std_logic_vector ( 22 downto 0 ) := "00111111000000011110100";

Signal ProductNode_POSIT1791Output_2215: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1793weight : std_logic_vector ( 22 downto 0 ) := "00111111101111110000101";

Signal ProductNode_POSIT1793Output_2217: std_logic_vector (22 downto 0);
Signal SumNode_POSIT424Output_2218: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1794Output_2219: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1799weight : std_logic_vector ( 22 downto 0 ) := "00111111000000011110100";

Signal ProductNode_POSIT1799Output_2225: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1801weight : std_logic_vector ( 22 downto 0 ) := "00111111101111110000101";

Signal ProductNode_POSIT1801Output_2227: std_logic_vector (22 downto 0);
Signal SumNode_POSIT426Output_2228: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1802Output_2229: std_logic_vector (22 downto 0);
Signal SumNode_POSIT427Output_2230: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1803Output_2231: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1809weight : std_logic_vector ( 22 downto 0 ) := "00111110001111100011101";

Signal ProductNode_POSIT1809Output_2238: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1811weight : std_logic_vector ( 22 downto 0 ) := "00111111111010000011100";

Signal ProductNode_POSIT1811Output_2240: std_logic_vector (22 downto 0);
Signal SumNode_POSIT429Output_2241: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1812Output_2242: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1817weight : std_logic_vector ( 22 downto 0 ) := "00111110001111100011101";

Signal ProductNode_POSIT1817Output_2248: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1819weight : std_logic_vector ( 22 downto 0 ) := "00111111111010000011100";

Signal ProductNode_POSIT1819Output_2250: std_logic_vector (22 downto 0);
Signal SumNode_POSIT431Output_2251: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1820Output_2252: std_logic_vector (22 downto 0);
Signal SumNode_POSIT432Output_2253: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1821Output_2254: std_logic_vector (22 downto 0);
Signal SumNode_POSIT433Output_2255: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1822Output_2256: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1849weight : std_logic_vector ( 22 downto 0 ) := "00111111111111100101101";

Signal ProductNode_POSIT1849Output_2287: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1853weight : std_logic_vector ( 22 downto 0 ) := "00111100010100101001100";

Signal ProductNode_POSIT1853Output_2292: std_logic_vector (22 downto 0);
Signal SumNode_POSIT439Output_2293: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1854Output_2294: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1881weight : std_logic_vector ( 22 downto 0 ) := "00111111111111111101111";

Signal ProductNode_POSIT1881Output_2325: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1885weight : std_logic_vector ( 22 downto 0 ) := "00111010100001000001111";

Signal ProductNode_POSIT1885Output_2330: std_logic_vector (22 downto 0);
Signal SumNode_POSIT445Output_2331: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1886Output_2332: std_logic_vector (22 downto 0);
Signal SumNode_POSIT446Output_2333: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1887Output_2334: std_logic_vector (22 downto 0);
Signal SumNode_POSIT447Output_2335: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1888Output_2336: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1890weight : std_logic_vector ( 22 downto 0 ) := "00111111011011011100000";

Signal ProductNode_POSIT1890Output_2338: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1927Output_2386: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1951weight : std_logic_vector ( 22 downto 0 ) := "00111110000110100001001";

Signal ProductNode_POSIT1951Output_2413: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1952weight : std_logic_vector ( 22 downto 0 ) := "00111111111011001011110";

Signal ProductNode_POSIT1952Output_2414: std_logic_vector (22 downto 0);
Signal SumNode_POSIT462Output_2415: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1953Output_2416: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1954weight : std_logic_vector ( 22 downto 0 ) := "00111111111001011010011";

Signal ProductNode_POSIT1954Output_2417: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1955weight : std_logic_vector ( 22 downto 0 ) := "00111001111101100110101";

Signal ProductNode_POSIT1955Output_2418: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1956weight : std_logic_vector ( 22 downto 0 ) := "00111111111111111111000";

Signal ProductNode_POSIT1956Output_2419: std_logic_vector (22 downto 0);
Signal SumNode_POSIT463Output_2420: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1957Output_2421: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1958weight : std_logic_vector ( 22 downto 0 ) := "00111110010100101100100";

Signal ProductNode_POSIT1958Output_2422: std_logic_vector (22 downto 0);
Signal SumNode_POSIT464Output_2423: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1959Output_2424: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1986weight : std_logic_vector ( 22 downto 0 ) := "00111111110100111101100";

Signal ProductNode_POSIT1986Output_2455: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1990weight : std_logic_vector ( 22 downto 0 ) := "00111110101100001001110";

Signal ProductNode_POSIT1990Output_2460: std_logic_vector (22 downto 0);
Signal SumNode_POSIT470Output_2461: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1991Output_2462: std_logic_vector (22 downto 0);
Signal SumNode_POSIT471Output_2463: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1992Output_2464: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT1994weight : std_logic_vector ( 22 downto 0 ) := "00111111101101111001001";

Signal ProductNode_POSIT1994Output_2466: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2031Output_2514: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2058weight : std_logic_vector ( 22 downto 0 ) := "00111111110010101000000";

Signal ProductNode_POSIT2058Output_2545: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2062weight : std_logic_vector ( 22 downto 0 ) := "00111110110101011111111";

Signal ProductNode_POSIT2062Output_2550: std_logic_vector (22 downto 0);
Signal SumNode_POSIT488Output_2551: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2063Output_2552: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2090weight : std_logic_vector ( 22 downto 0 ) := "00111111101101101101100";

Signal ProductNode_POSIT2090Output_2583: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2094weight : std_logic_vector ( 22 downto 0 ) := "00111111000100100100111";

Signal ProductNode_POSIT2094Output_2588: std_logic_vector (22 downto 0);
Signal SumNode_POSIT494Output_2589: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2095Output_2590: std_logic_vector (22 downto 0);
Signal SumNode_POSIT495Output_2591: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2096Output_2592: std_logic_vector (22 downto 0);
Signal SumNode_POSIT496Output_2593: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2097Output_2594: std_logic_vector (22 downto 0);
Signal SumNode_POSIT497Output_2595: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2098Output_2596: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2101weight : std_logic_vector ( 22 downto 0 ) := "00111110011000001010100";

Signal ProductNode_POSIT2101Output_2599: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2118Output_2621: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2119weight : std_logic_vector ( 22 downto 0 ) := "00111111111000111110101";

Signal ProductNode_POSIT2119Output_2622: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2136Output_2644: std_logic_vector (22 downto 0);
Signal SumNode_POSIT508Output_2645: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2137Output_2646: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2164weight : std_logic_vector ( 22 downto 0 ) := "00111111111110000111011";

Signal ProductNode_POSIT2164Output_2677: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2168weight : std_logic_vector ( 22 downto 0 ) := "00111101011100010001110";

Signal ProductNode_POSIT2168Output_2682: std_logic_vector (22 downto 0);
Signal SumNode_POSIT514Output_2683: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2169Output_2684: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2196weight : std_logic_vector ( 22 downto 0 ) := "00111111111010100100111";

Signal ProductNode_POSIT2196Output_2715: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2200weight : std_logic_vector ( 22 downto 0 ) := "00111110001011011000011";

Signal ProductNode_POSIT2200Output_2720: std_logic_vector (22 downto 0);
Signal SumNode_POSIT520Output_2721: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2201Output_2722: std_logic_vector (22 downto 0);
Signal SumNode_POSIT521Output_2723: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2202Output_2724: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2222Output_2749: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2240Output_2772: std_logic_vector (22 downto 0);
Signal SumNode_POSIT532Output_2773: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2241Output_2774: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2268weight : std_logic_vector ( 22 downto 0 ) := "00111111110101101110000";

Signal ProductNode_POSIT2268Output_2805: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2272weight : std_logic_vector ( 22 downto 0 ) := "00111110101001000111101";

Signal ProductNode_POSIT2272Output_2810: std_logic_vector (22 downto 0);
Signal SumNode_POSIT538Output_2811: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2273Output_2812: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2300weight : std_logic_vector ( 22 downto 0 ) := "00111111111000011101001";

Signal ProductNode_POSIT2300Output_2843: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2304weight : std_logic_vector ( 22 downto 0 ) := "00111110011100010110101";

Signal ProductNode_POSIT2304Output_2848: std_logic_vector (22 downto 0);
Signal SumNode_POSIT544Output_2849: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2305Output_2850: std_logic_vector (22 downto 0);
Signal SumNode_POSIT545Output_2851: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2306Output_2852: std_logic_vector (22 downto 0);
Signal SumNode_POSIT546Output_2853: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2307Output_2854: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2346Output_2904: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2373weight : std_logic_vector ( 22 downto 0 ) := "00111111110010101111110";

Signal ProductNode_POSIT2373Output_2935: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2377weight : std_logic_vector ( 22 downto 0 ) := "00111110110101000000100";

Signal ProductNode_POSIT2377Output_2940: std_logic_vector (22 downto 0);
Signal SumNode_POSIT563Output_2941: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2378Output_2942: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2405weight : std_logic_vector ( 22 downto 0 ) := "00111111101100011011010";

Signal ProductNode_POSIT2405Output_2973: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2409weight : std_logic_vector ( 22 downto 0 ) := "00111111000111001001011";

Signal ProductNode_POSIT2409Output_2978: std_logic_vector (22 downto 0);
Signal SumNode_POSIT569Output_2979: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2410Output_2980: std_logic_vector (22 downto 0);
Signal SumNode_POSIT570Output_2981: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2411Output_2982: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2450Output_3032: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2477weight : std_logic_vector ( 22 downto 0 ) := "00111111101100100011100";

Signal ProductNode_POSIT2477Output_3063: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2481weight : std_logic_vector ( 22 downto 0 ) := "00111111000110111000110";

Signal ProductNode_POSIT2481Output_3068: std_logic_vector (22 downto 0);
Signal SumNode_POSIT587Output_3069: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2482Output_3070: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2509weight : std_logic_vector ( 22 downto 0 ) := "00111111100001101001010";

Signal ProductNode_POSIT2509Output_3101: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2513weight : std_logic_vector ( 22 downto 0 ) := "00111111011100101101011";

Signal ProductNode_POSIT2513Output_3106: std_logic_vector (22 downto 0);
Signal SumNode_POSIT593Output_3107: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2514Output_3108: std_logic_vector (22 downto 0);
Signal SumNode_POSIT594Output_3109: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2515Output_3110: std_logic_vector (22 downto 0);
Signal SumNode_POSIT595Output_3111: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2516Output_3112: std_logic_vector (22 downto 0);
Signal SumNode_POSIT596Output_3113: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2517Output_3114: std_logic_vector (22 downto 0);
Signal SumNode_POSIT597Output_3115: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2518Output_3116: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2519weight : std_logic_vector ( 22 downto 0 ) := "00111111101011110001010";

Signal ProductNode_POSIT2519Output_3117: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2520weight : std_logic_vector ( 22 downto 0 ) := "00111111100010010001111";

Signal ProductNode_POSIT2520Output_3118: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2521weight : std_logic_vector ( 22 downto 0 ) := "00111110010011011101101";

Signal ProductNode_POSIT2521Output_3119: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2522weight : std_logic_vector ( 22 downto 0 ) := "00111110000100110001000";

Signal ProductNode_POSIT2522Output_3120: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2523weight : std_logic_vector ( 22 downto 0 ) := "00111111111011011001110";

Signal ProductNode_POSIT2523Output_3121: std_logic_vector (22 downto 0);
Signal SumNode_POSIT598Output_3122: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2524Output_3123: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2529Output_3129: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2530weight : std_logic_vector ( 22 downto 0 ) := "00111100101110010011110";

Signal ProductNode_POSIT2530Output_3130: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2531weight : std_logic_vector ( 22 downto 0 ) := "00111111111111010001101";

Signal ProductNode_POSIT2531Output_3131: std_logic_vector (22 downto 0);
Signal SumNode_POSIT600Output_3132: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2532Output_3133: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2537Output_3139: std_logic_vector (22 downto 0);
Signal SumNode_POSIT602Output_3140: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2538Output_3141: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2539weight : std_logic_vector ( 22 downto 0 ) := "00111111111001100100010";

Signal ProductNode_POSIT2539Output_3142: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2547Output_3152: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2555Output_3162: std_logic_vector (22 downto 0);
Signal SumNode_POSIT607Output_3163: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2556Output_3164: std_logic_vector (22 downto 0);
Signal SumNode_POSIT608Output_3165: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2557Output_3166: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2581weight : std_logic_vector ( 22 downto 0 ) := "00111110101011100011000";

Signal ProductNode_POSIT2581Output_3193: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2582weight : std_logic_vector ( 22 downto 0 ) := "00111111110101000111001";

Signal ProductNode_POSIT2582Output_3194: std_logic_vector (22 downto 0);
Signal SumNode_POSIT612Output_3195: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2583Output_3196: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2584weight : std_logic_vector ( 22 downto 0 ) := "00111111111111100101100";

Signal ProductNode_POSIT2584Output_3197: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2585weight : std_logic_vector ( 22 downto 0 ) := "00111100110100000110111";

Signal ProductNode_POSIT2585Output_3198: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2586weight : std_logic_vector ( 22 downto 0 ) := "00111111111111001011111";

Signal ProductNode_POSIT2586Output_3199: std_logic_vector (22 downto 0);
Signal SumNode_POSIT613Output_3200: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2587Output_3201: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2588weight : std_logic_vector ( 22 downto 0 ) := "00111100010100111011011";

Signal ProductNode_POSIT2588Output_3202: std_logic_vector (22 downto 0);
Signal SumNode_POSIT614Output_3203: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2589Output_3204: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2616weight : std_logic_vector ( 22 downto 0 ) := "00111111111110010011111";

Signal ProductNode_POSIT2616Output_3235: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2620weight : std_logic_vector ( 22 downto 0 ) := "00111101010110000001110";

Signal ProductNode_POSIT2620Output_3240: std_logic_vector (22 downto 0);
Signal SumNode_POSIT620Output_3241: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2621Output_3242: std_logic_vector (22 downto 0);
Signal SumNode_POSIT621Output_3243: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2622Output_3244: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2623weight : std_logic_vector ( 22 downto 0 ) := "00111111111110100010010";

Signal ProductNode_POSIT2623Output_3245: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2624weight : std_logic_vector ( 22 downto 0 ) := "00111111000100001101101";

Signal ProductNode_POSIT2624Output_3246: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2633Output_3257: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2641Output_3267: std_logic_vector (22 downto 0);
Signal SumNode_POSIT626Output_3268: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2642Output_3269: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2651Output_3280: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2659Output_3290: std_logic_vector (22 downto 0);
Signal SumNode_POSIT631Output_3291: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2660Output_3292: std_logic_vector (22 downto 0);
Signal SumNode_POSIT632Output_3293: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2661Output_3294: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2688weight : std_logic_vector ( 22 downto 0 ) := "00111111111111100101101";

Signal ProductNode_POSIT2688Output_3325: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2692weight : std_logic_vector ( 22 downto 0 ) := "00111100010100101001100";

Signal ProductNode_POSIT2692Output_3330: std_logic_vector (22 downto 0);
Signal SumNode_POSIT638Output_3331: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2693Output_3332: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2720weight : std_logic_vector ( 22 downto 0 ) := "00111111111111111101111";

Signal ProductNode_POSIT2720Output_3363: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2724weight : std_logic_vector ( 22 downto 0 ) := "00111010100001000001111";

Signal ProductNode_POSIT2724Output_3368: std_logic_vector (22 downto 0);
Signal SumNode_POSIT644Output_3369: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2725Output_3370: std_logic_vector (22 downto 0);
Signal SumNode_POSIT645Output_3371: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2726Output_3372: std_logic_vector (22 downto 0);
Signal SumNode_POSIT646Output_3373: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2727Output_3374: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2729weight : std_logic_vector ( 22 downto 0 ) := "00111111011011011100000";

Signal ProductNode_POSIT2729Output_3376: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2766Output_3424: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2790weight : std_logic_vector ( 22 downto 0 ) := "00111101010000011111101";

Signal ProductNode_POSIT2790Output_3451: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2791weight : std_logic_vector ( 22 downto 0 ) := "00111111111110011111000";

Signal ProductNode_POSIT2791Output_3452: std_logic_vector (22 downto 0);
Signal SumNode_POSIT661Output_3453: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2792Output_3454: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2793weight : std_logic_vector ( 22 downto 0 ) := "00111111111001011010011";

Signal ProductNode_POSIT2793Output_3455: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2794weight : std_logic_vector ( 22 downto 0 ) := "00110111010010010101001";

Signal ProductNode_POSIT2794Output_3456: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2795weight : std_logic_vector ( 22 downto 0 ) := "00111111111111111111111";

Signal ProductNode_POSIT2795Output_3457: std_logic_vector (22 downto 0);
Signal SumNode_POSIT662Output_3458: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2796Output_3459: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2797weight : std_logic_vector ( 22 downto 0 ) := "00111110010100101100100";

Signal ProductNode_POSIT2797Output_3460: std_logic_vector (22 downto 0);
Signal SumNode_POSIT663Output_3461: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2798Output_3462: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2825weight : std_logic_vector ( 22 downto 0 ) := "00111111110100111101100";

Signal ProductNode_POSIT2825Output_3493: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2829weight : std_logic_vector ( 22 downto 0 ) := "00111110101100001001110";

Signal ProductNode_POSIT2829Output_3498: std_logic_vector (22 downto 0);
Signal SumNode_POSIT669Output_3499: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2830Output_3500: std_logic_vector (22 downto 0);
Signal SumNode_POSIT670Output_3501: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2831Output_3502: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2833weight : std_logic_vector ( 22 downto 0 ) := "00111111101101111001001";

Signal ProductNode_POSIT2833Output_3504: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2870Output_3552: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2897weight : std_logic_vector ( 22 downto 0 ) := "00111111110010101000000";

Signal ProductNode_POSIT2897Output_3583: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2901weight : std_logic_vector ( 22 downto 0 ) := "00111110110101011111111";

Signal ProductNode_POSIT2901Output_3588: std_logic_vector (22 downto 0);
Signal SumNode_POSIT687Output_3589: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2902Output_3590: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2929weight : std_logic_vector ( 22 downto 0 ) := "00111111101101101101100";

Signal ProductNode_POSIT2929Output_3621: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2933weight : std_logic_vector ( 22 downto 0 ) := "00111111000100100100111";

Signal ProductNode_POSIT2933Output_3626: std_logic_vector (22 downto 0);
Signal SumNode_POSIT693Output_3627: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2934Output_3628: std_logic_vector (22 downto 0);
Signal SumNode_POSIT694Output_3629: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2935Output_3630: std_logic_vector (22 downto 0);
Signal SumNode_POSIT695Output_3631: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2936Output_3632: std_logic_vector (22 downto 0);
Signal SumNode_POSIT696Output_3633: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2937Output_3634: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2940weight : std_logic_vector ( 22 downto 0 ) := "00111101111001011101111";

Signal ProductNode_POSIT2940Output_3637: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2957Output_3659: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2958weight : std_logic_vector ( 22 downto 0 ) := "00111111111100011010001";

Signal ProductNode_POSIT2958Output_3660: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2975Output_3682: std_logic_vector (22 downto 0);
Signal SumNode_POSIT707Output_3683: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT2976Output_3684: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3003weight : std_logic_vector ( 22 downto 0 ) := "00111111111110000111011";

Signal ProductNode_POSIT3003Output_3715: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3007weight : std_logic_vector ( 22 downto 0 ) := "00111101011100010001110";

Signal ProductNode_POSIT3007Output_3720: std_logic_vector (22 downto 0);
Signal SumNode_POSIT713Output_3721: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3008Output_3722: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3035weight : std_logic_vector ( 22 downto 0 ) := "00111111111010100100111";

Signal ProductNode_POSIT3035Output_3753: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3039weight : std_logic_vector ( 22 downto 0 ) := "00111110001011011000011";

Signal ProductNode_POSIT3039Output_3758: std_logic_vector (22 downto 0);
Signal SumNode_POSIT719Output_3759: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3040Output_3760: std_logic_vector (22 downto 0);
Signal SumNode_POSIT720Output_3761: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3041Output_3762: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3061Output_3787: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3079Output_3810: std_logic_vector (22 downto 0);
Signal SumNode_POSIT731Output_3811: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3080Output_3812: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3107weight : std_logic_vector ( 22 downto 0 ) := "00111111110101101110000";

Signal ProductNode_POSIT3107Output_3843: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3111weight : std_logic_vector ( 22 downto 0 ) := "00111110101001000111101";

Signal ProductNode_POSIT3111Output_3848: std_logic_vector (22 downto 0);
Signal SumNode_POSIT737Output_3849: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3112Output_3850: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3139weight : std_logic_vector ( 22 downto 0 ) := "00111111111000011101001";

Signal ProductNode_POSIT3139Output_3881: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3143weight : std_logic_vector ( 22 downto 0 ) := "00111110011100010110101";

Signal ProductNode_POSIT3143Output_3886: std_logic_vector (22 downto 0);
Signal SumNode_POSIT743Output_3887: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3144Output_3888: std_logic_vector (22 downto 0);
Signal SumNode_POSIT744Output_3889: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3145Output_3890: std_logic_vector (22 downto 0);
Signal SumNode_POSIT745Output_3891: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3146Output_3892: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3185Output_3942: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3212weight : std_logic_vector ( 22 downto 0 ) := "00111111110010101111110";

Signal ProductNode_POSIT3212Output_3973: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3216weight : std_logic_vector ( 22 downto 0 ) := "00111110110101000000100";

Signal ProductNode_POSIT3216Output_3978: std_logic_vector (22 downto 0);
Signal SumNode_POSIT762Output_3979: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3217Output_3980: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3244weight : std_logic_vector ( 22 downto 0 ) := "00111111101100011011010";

Signal ProductNode_POSIT3244Output_4011: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3248weight : std_logic_vector ( 22 downto 0 ) := "00111111000111001001011";

Signal ProductNode_POSIT3248Output_4016: std_logic_vector (22 downto 0);
Signal SumNode_POSIT768Output_4017: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3249Output_4018: std_logic_vector (22 downto 0);
Signal SumNode_POSIT769Output_4019: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3250Output_4020: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3289Output_4070: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3316weight : std_logic_vector ( 22 downto 0 ) := "00111111101100100011100";

Signal ProductNode_POSIT3316Output_4101: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3320weight : std_logic_vector ( 22 downto 0 ) := "00111111000110111000110";

Signal ProductNode_POSIT3320Output_4106: std_logic_vector (22 downto 0);
Signal SumNode_POSIT786Output_4107: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3321Output_4108: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3348weight : std_logic_vector ( 22 downto 0 ) := "00111111100001101001010";

Signal ProductNode_POSIT3348Output_4139: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3352weight : std_logic_vector ( 22 downto 0 ) := "00111111011100101101011";

Signal ProductNode_POSIT3352Output_4144: std_logic_vector (22 downto 0);
Signal SumNode_POSIT792Output_4145: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3353Output_4146: std_logic_vector (22 downto 0);
Signal SumNode_POSIT793Output_4147: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3354Output_4148: std_logic_vector (22 downto 0);
Signal SumNode_POSIT794Output_4149: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3355Output_4150: std_logic_vector (22 downto 0);
Signal SumNode_POSIT795Output_4151: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3356Output_4152: std_logic_vector (22 downto 0);
Signal SumNode_POSIT796Output_4153: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3357Output_4154: std_logic_vector (22 downto 0);
Signal SumNode_POSIT797Output_4155: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3358Output_4156: std_logic_vector (22 downto 0);
Signal SumNode_POSIT798Output_4157: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3359Output_4158: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3361weight : std_logic_vector ( 22 downto 0 ) := "00111111110100101110111";

Signal ProductNode_POSIT3361Output_4160: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3363weight : std_logic_vector ( 22 downto 0 ) := "00111110110110110001010";

Signal ProductNode_POSIT3363Output_4162: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3364weight : std_logic_vector ( 22 downto 0 ) := "00111111110010010011101";

Signal ProductNode_POSIT3364Output_4163: std_logic_vector (22 downto 0);
Signal SumNode_POSIT799Output_4164: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3365Output_4165: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3370Output_4171: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3371weight : std_logic_vector ( 22 downto 0 ) := "00111110100101111111111";

Signal ProductNode_POSIT3371Output_4172: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3372weight : std_logic_vector ( 22 downto 0 ) := "00111111110110100000000";

Signal ProductNode_POSIT3372Output_4173: std_logic_vector (22 downto 0);
Signal SumNode_POSIT801Output_4174: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3373Output_4175: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3378Output_4181: std_logic_vector (22 downto 0);
Signal SumNode_POSIT803Output_4182: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3379Output_4183: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3388Output_4194: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3396Output_4204: std_logic_vector (22 downto 0);
Signal SumNode_POSIT808Output_4205: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3397Output_4206: std_logic_vector (22 downto 0);
Signal SumNode_POSIT809Output_4207: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3398Output_4208: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3401weight : std_logic_vector ( 22 downto 0 ) := "00111111010000010010011";

Signal ProductNode_POSIT3401Output_4211: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3402weight : std_logic_vector ( 22 downto 0 ) := "00111111000011010101101";

Signal ProductNode_POSIT3402Output_4212: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3403weight : std_logic_vector ( 22 downto 0 ) := "00111111110010101100001";

Signal ProductNode_POSIT3403Output_4213: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3405weight : std_logic_vector ( 22 downto 0 ) := "00111111111010111011100";

Signal ProductNode_POSIT3405Output_4215: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3406weight : std_logic_vector ( 22 downto 0 ) := "00111110011010010100011";

Signal ProductNode_POSIT3406Output_4216: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3407weight : std_logic_vector ( 22 downto 0 ) := "00111111101101100111110";

Signal ProductNode_POSIT3407Output_4217: std_logic_vector (22 downto 0);
Signal SumNode_POSIT810Output_4218: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3408Output_4219: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3409weight : std_logic_vector ( 22 downto 0 ) := "00111111000011101010101";

Signal ProductNode_POSIT3409Output_4220: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3412weight : std_logic_vector ( 22 downto 0 ) := "00111111101110010101001";

Signal ProductNode_POSIT3412Output_4223: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3413weight : std_logic_vector ( 22 downto 0 ) := "00111111011001101110010";

Signal ProductNode_POSIT3413Output_4224: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3416weight : std_logic_vector ( 22 downto 0 ) := "00111111111000101101011";

Signal ProductNode_POSIT3416Output_4227: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3417weight : std_logic_vector ( 22 downto 0 ) := "00111111001101100010000";

Signal ProductNode_POSIT3417Output_4228: std_logic_vector (22 downto 0);
Signal SumNode_POSIT811Output_4229: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3418Output_4230: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3419weight : std_logic_vector ( 22 downto 0 ) := "00111110100000010010111";

Signal ProductNode_POSIT3419Output_4231: std_logic_vector (22 downto 0);
Signal SumNode_POSIT812Output_4232: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3420Output_4233: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3421weight : std_logic_vector ( 22 downto 0 ) := "00111111111000110110110";

Signal ProductNode_POSIT3421Output_4234: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3430Output_4246: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3433weight : std_logic_vector ( 22 downto 0 ) := "00111111001010011111000";

Signal ProductNode_POSIT3433Output_4249: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3434weight : std_logic_vector ( 22 downto 0 ) := "00111110111001100001111";

Signal ProductNode_POSIT3434Output_4250: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3435weight : std_logic_vector ( 22 downto 0 ) := "00111111110000011101000";

Signal ProductNode_POSIT3435Output_4251: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3437weight : std_logic_vector ( 22 downto 0 ) := "00111111111110110011010";

Signal ProductNode_POSIT3437Output_4253: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3438weight : std_logic_vector ( 22 downto 0 ) := "00111101100000000101110";

Signal ProductNode_POSIT3438Output_4254: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3439weight : std_logic_vector ( 22 downto 0 ) := "00111111100101000110011";

Signal ProductNode_POSIT3439Output_4255: std_logic_vector (22 downto 0);
Signal SumNode_POSIT816Output_4256: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3440Output_4257: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3441weight : std_logic_vector ( 22 downto 0 ) := "00111111000011101010101";

Signal ProductNode_POSIT3441Output_4258: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3444weight : std_logic_vector ( 22 downto 0 ) := "00111111110001100111100";

Signal ProductNode_POSIT3444Output_4261: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3445weight : std_logic_vector ( 22 downto 0 ) := "00111111010101111001100";

Signal ProductNode_POSIT3445Output_4262: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3448weight : std_logic_vector ( 22 downto 0 ) := "00111111111101111111101";

Signal ProductNode_POSIT3448Output_4265: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3449weight : std_logic_vector ( 22 downto 0 ) := "00111110100010110011010";

Signal ProductNode_POSIT3449Output_4266: std_logic_vector (22 downto 0);
Signal SumNode_POSIT817Output_4267: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3450Output_4268: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3451weight : std_logic_vector ( 22 downto 0 ) := "00111110100000010010111";

Signal ProductNode_POSIT3451Output_4269: std_logic_vector (22 downto 0);
Signal SumNode_POSIT818Output_4270: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3452Output_4271: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3453weight : std_logic_vector ( 22 downto 0 ) := "00111111101100111001011";

Signal ProductNode_POSIT3453Output_4272: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3462Output_4284: std_logic_vector (22 downto 0);
Signal SumNode_POSIT822Output_4285: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3463Output_4286: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3465weight : std_logic_vector ( 22 downto 0 ) := "00111111100010110101010";

Signal ProductNode_POSIT3465Output_4288: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3474Output_4299: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3482Output_4309: std_logic_vector (22 downto 0);
Signal SumNode_POSIT827Output_4310: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3483Output_4311: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3492Output_4322: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3500Output_4332: std_logic_vector (22 downto 0);
Signal SumNode_POSIT832Output_4333: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3501Output_4334: std_logic_vector (22 downto 0);
Signal SumNode_POSIT833Output_4335: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3502Output_4336: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3525weight : std_logic_vector ( 22 downto 0 ) := "00111110011001001001101";

Signal ProductNode_POSIT3525Output_4362: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3534Output_4374: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3557weight : std_logic_vector ( 22 downto 0 ) := "00111111000110001101000";

Signal ProductNode_POSIT3557Output_4400: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3566Output_4412: std_logic_vector (22 downto 0);
Signal SumNode_POSIT846Output_4413: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3567Output_4414: std_logic_vector (22 downto 0);
Signal SumNode_POSIT847Output_4415: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3568Output_4416: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3570weight : std_logic_vector ( 22 downto 0 ) := "00111110101101000100010";

Signal ProductNode_POSIT3570Output_4418: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3607Output_4466: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3639Output_4504: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3671Output_4542: std_logic_vector (22 downto 0);
Signal SumNode_POSIT871Output_4543: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3672Output_4544: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3674weight : std_logic_vector ( 22 downto 0 ) := "00111111011010010101010";

Signal ProductNode_POSIT3674Output_4546: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3711Output_4594: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3743Output_4632: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3775Output_4670: std_logic_vector (22 downto 0);
Signal SumNode_POSIT895Output_4671: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3776Output_4672: std_logic_vector (22 downto 0);
Signal SumNode_POSIT896Output_4673: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3777Output_4674: std_logic_vector (22 downto 0);
Signal SumNode_POSIT897Output_4675: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3778Output_4676: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3798Output_4701: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3816Output_4724: std_logic_vector (22 downto 0);
Signal SumNode_POSIT908Output_4725: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3817Output_4726: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3822weight : std_logic_vector ( 22 downto 0 ) := "00111110110101001111010";

Signal ProductNode_POSIT3822Output_4731: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3826weight : std_logic_vector ( 22 downto 0 ) := "00111111000100110000010";

Signal ProductNode_POSIT3826Output_4735: std_logic_vector (22 downto 0);
Signal SumNode_POSIT909Output_4736: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3827Output_4737: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3828weight : std_logic_vector ( 22 downto 0 ) := "00111110001101100110000";

Signal ProductNode_POSIT3828Output_4738: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3832weight : std_logic_vector ( 22 downto 0 ) := "00111111100011001000110";

Signal ProductNode_POSIT3832Output_4742: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3836weight : std_logic_vector ( 22 downto 0 ) := "00111111101001001110111";

Signal ProductNode_POSIT3836Output_4746: std_logic_vector (22 downto 0);
Signal SumNode_POSIT910Output_4747: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3837Output_4748: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3838weight : std_logic_vector ( 22 downto 0 ) := "00111101001100001111101";

Signal ProductNode_POSIT3838Output_4749: std_logic_vector (22 downto 0);
Signal SumNode_POSIT911Output_4750: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3839Output_4751: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3840weight : std_logic_vector ( 22 downto 0 ) := "00111111101111011010100";

Signal ProductNode_POSIT3840Output_4752: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3849Output_4764: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3854weight : std_logic_vector ( 22 downto 0 ) := "00111110111110001011110";

Signal ProductNode_POSIT3854Output_4769: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3858weight : std_logic_vector ( 22 downto 0 ) := "00111111010101110011001";

Signal ProductNode_POSIT3858Output_4773: std_logic_vector (22 downto 0);
Signal SumNode_POSIT915Output_4774: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3859Output_4775: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3860weight : std_logic_vector ( 22 downto 0 ) := "00111110001101100110000";

Signal ProductNode_POSIT3860Output_4776: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3864weight : std_logic_vector ( 22 downto 0 ) := "00111111100101000011001";

Signal ProductNode_POSIT3864Output_4780: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3868weight : std_logic_vector ( 22 downto 0 ) := "00111111110111010011001";

Signal ProductNode_POSIT3868Output_4784: std_logic_vector (22 downto 0);
Signal SumNode_POSIT916Output_4785: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3869Output_4786: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3870weight : std_logic_vector ( 22 downto 0 ) := "00111101001100001111101";

Signal ProductNode_POSIT3870Output_4787: std_logic_vector (22 downto 0);
Signal SumNode_POSIT917Output_4788: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3871Output_4789: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3872weight : std_logic_vector ( 22 downto 0 ) := "00111111100101000101011";

Signal ProductNode_POSIT3872Output_4790: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3881Output_4802: std_logic_vector (22 downto 0);
Signal SumNode_POSIT921Output_4803: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3882Output_4804: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3902Output_4829: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3920Output_4852: std_logic_vector (22 downto 0);
Signal SumNode_POSIT932Output_4853: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3921Output_4854: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3944weight : std_logic_vector ( 22 downto 0 ) := "00111111000001001010110";

Signal ProductNode_POSIT3944Output_4880: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3953Output_4892: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3976weight : std_logic_vector ( 22 downto 0 ) := "00111111010101110101001";

Signal ProductNode_POSIT3976Output_4918: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3985Output_4930: std_logic_vector (22 downto 0);
Signal SumNode_POSIT945Output_4931: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3986Output_4932: std_logic_vector (22 downto 0);
Signal SumNode_POSIT946Output_4933: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT3987Output_4934: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4026Output_4984: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4058Output_5022: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4090Output_5060: std_logic_vector (22 downto 0);
Signal SumNode_POSIT970Output_5061: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4091Output_5062: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4130Output_5112: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4162Output_5150: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4194Output_5188: std_logic_vector (22 downto 0);
Signal SumNode_POSIT994Output_5189: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4195Output_5190: std_logic_vector (22 downto 0);
Signal SumNode_POSIT995Output_5191: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4196Output_5192: std_logic_vector (22 downto 0);
Signal SumNode_POSIT996Output_5193: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4197Output_5194: std_logic_vector (22 downto 0);
Signal SumNode_POSIT997Output_5195: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4198Output_5196: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4200weight : std_logic_vector ( 22 downto 0 ) := "00111111110100101110111";

Signal ProductNode_POSIT4200Output_5198: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4202weight : std_logic_vector ( 22 downto 0 ) := "00111110000001100101101";

Signal ProductNode_POSIT4202Output_5200: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4203weight : std_logic_vector ( 22 downto 0 ) := "00111111111011110011010";

Signal ProductNode_POSIT4203Output_5201: std_logic_vector (22 downto 0);
Signal SumNode_POSIT998Output_5202: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4204Output_5203: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4209Output_5209: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4210weight : std_logic_vector ( 22 downto 0 ) := "00111101010111111111000";

Signal ProductNode_POSIT4210Output_5210: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4211weight : std_logic_vector ( 22 downto 0 ) := "00111111111110010000000";

Signal ProductNode_POSIT4211Output_5211: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1000Output_5212: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4212Output_5213: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4217Output_5219: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1002Output_5220: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4218Output_5221: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4227Output_5232: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4235Output_5242: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1007Output_5243: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4236Output_5244: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1008Output_5245: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4237Output_5246: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4248weight : std_logic_vector ( 22 downto 0 ) := "00111111101110001010101";

Signal ProductNode_POSIT4248Output_5258: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4258weight : std_logic_vector ( 22 downto 0 ) := "00111111110111111011010";

Signal ProductNode_POSIT4258Output_5269: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1011Output_5270: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4259Output_5271: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4260weight : std_logic_vector ( 22 downto 0 ) := "00111111111000110110110";

Signal ProductNode_POSIT4260Output_5272: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4269Output_5284: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4280weight : std_logic_vector ( 22 downto 0 ) := "00111111101110001010101";

Signal ProductNode_POSIT4280Output_5296: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4290weight : std_logic_vector ( 22 downto 0 ) := "00111111110111111011010";

Signal ProductNode_POSIT4290Output_5307: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1017Output_5308: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4291Output_5309: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4292weight : std_logic_vector ( 22 downto 0 ) := "00111111101100111001011";

Signal ProductNode_POSIT4292Output_5310: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4301Output_5322: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1021Output_5323: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4302Output_5324: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4304weight : std_logic_vector ( 22 downto 0 ) := "00111111100010110101010";

Signal ProductNode_POSIT4304Output_5326: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4313Output_5337: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4321Output_5347: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1026Output_5348: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4322Output_5349: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4331Output_5360: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4339Output_5370: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1031Output_5371: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4340Output_5372: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1032Output_5373: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4341Output_5374: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4364weight : std_logic_vector ( 22 downto 0 ) := "00111110011001001001101";

Signal ProductNode_POSIT4364Output_5400: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4373Output_5412: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4396weight : std_logic_vector ( 22 downto 0 ) := "00111111000110001101000";

Signal ProductNode_POSIT4396Output_5438: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4405Output_5450: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1045Output_5451: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4406Output_5452: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1046Output_5453: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4407Output_5454: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4409weight : std_logic_vector ( 22 downto 0 ) := "00111110101101000100010";

Signal ProductNode_POSIT4409Output_5456: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4446Output_5504: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4478Output_5542: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4510Output_5580: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1070Output_5581: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4511Output_5582: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4513weight : std_logic_vector ( 22 downto 0 ) := "00111111011010010101010";

Signal ProductNode_POSIT4513Output_5584: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4550Output_5632: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4582Output_5670: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4614Output_5708: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1094Output_5709: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4615Output_5710: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1095Output_5711: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4616Output_5712: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1096Output_5713: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4617Output_5714: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4637Output_5739: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4655Output_5762: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1107Output_5763: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4656Output_5764: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4667weight : std_logic_vector ( 22 downto 0 ) := "00111111111010010011001";

Signal ProductNode_POSIT4667Output_5776: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4677weight : std_logic_vector ( 22 downto 0 ) := "00111111111110100111100";

Signal ProductNode_POSIT4677Output_5787: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1110Output_5788: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4678Output_5789: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4679weight : std_logic_vector ( 22 downto 0 ) := "00111111101111011010100";

Signal ProductNode_POSIT4679Output_5790: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4688Output_5802: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4699weight : std_logic_vector ( 22 downto 0 ) := "00111111111010010011001";

Signal ProductNode_POSIT4699Output_5814: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4709weight : std_logic_vector ( 22 downto 0 ) := "00111111111110100111100";

Signal ProductNode_POSIT4709Output_5825: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1116Output_5826: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4710Output_5827: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4711weight : std_logic_vector ( 22 downto 0 ) := "00111111100101000101011";

Signal ProductNode_POSIT4711Output_5828: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4720Output_5840: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1120Output_5841: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4721Output_5842: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4741Output_5867: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4759Output_5890: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1131Output_5891: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4760Output_5892: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4783weight : std_logic_vector ( 22 downto 0 ) := "00111111000001001010110";

Signal ProductNode_POSIT4783Output_5918: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4792Output_5930: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4815weight : std_logic_vector ( 22 downto 0 ) := "00111111010101110101001";

Signal ProductNode_POSIT4815Output_5956: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4824Output_5968: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1144Output_5969: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4825Output_5970: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1145Output_5971: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4826Output_5972: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4865Output_6022: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4897Output_6060: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4929Output_6098: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1169Output_6099: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4930Output_6100: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT4969Output_6150: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5001Output_6188: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5033Output_6226: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1193Output_6227: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5034Output_6228: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1194Output_6229: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5035Output_6230: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1195Output_6231: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5036Output_6232: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1196Output_6233: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5037Output_6234: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1197Output_6235: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5038Output_6236: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5040weight : std_logic_vector ( 22 downto 0 ) := "00111111001100010101001";

Signal ProductNode_POSIT5040Output_6238: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5042weight : std_logic_vector ( 22 downto 0 ) := "00111110010111101100001";

Signal ProductNode_POSIT5042Output_6240: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5043weight : std_logic_vector ( 22 downto 0 ) := "00111111111001000010011";

Signal ProductNode_POSIT5043Output_6241: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1198Output_6242: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5044Output_6243: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5049Output_6249: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5050weight : std_logic_vector ( 22 downto 0 ) := "00111101100010100110011";

Signal ProductNode_POSIT5050Output_6250: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5051weight : std_logic_vector ( 22 downto 0 ) := "00111111111101110101100";

Signal ProductNode_POSIT5051Output_6251: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1200Output_6252: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5052Output_6253: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5057Output_6259: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1202Output_6260: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5058Output_6261: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5067Output_6272: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5075Output_6282: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1207Output_6283: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5076Output_6284: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1208Output_6285: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5077Output_6286: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5109Output_6324: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5141Output_6362: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1221Output_6363: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5142Output_6364: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5144weight : std_logic_vector ( 22 downto 0 ) := "00111110100010010000110";

Signal ProductNode_POSIT5144Output_6366: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5153Output_6377: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5161Output_6387: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1226Output_6388: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5162Output_6389: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5171Output_6400: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5179Output_6410: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1231Output_6411: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5180Output_6412: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1232Output_6413: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5181Output_6414: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5213Output_6452: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5245Output_6490: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1245Output_6491: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5246Output_6492: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1246Output_6493: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5247Output_6494: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5249weight : std_logic_vector ( 22 downto 0 ) := "00111111101001110101011";

Signal ProductNode_POSIT5249Output_6496: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5286Output_6544: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5318Output_6582: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5350Output_6620: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1270Output_6621: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5351Output_6622: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5353weight : std_logic_vector ( 22 downto 0 ) := "00111111110111011011110";

Signal ProductNode_POSIT5353Output_6624: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5390Output_6672: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5422Output_6710: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5454Output_6748: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1294Output_6749: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5455Output_6750: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1295Output_6751: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5456Output_6752: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1296Output_6753: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5457Output_6754: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5477Output_6779: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5495Output_6802: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1307Output_6803: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5496Output_6804: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5528Output_6842: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5560Output_6880: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1320Output_6881: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5561Output_6882: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5581Output_6907: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5599Output_6930: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1331Output_6931: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5600Output_6932: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5632Output_6970: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5664Output_7008: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1344Output_7009: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5665Output_7010: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1345Output_7011: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5666Output_7012: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5705Output_7062: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5737Output_7100: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5769Output_7138: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1369Output_7139: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5770Output_7140: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5809Output_7190: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5841Output_7228: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5873Output_7266: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1393Output_7267: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5874Output_7268: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1394Output_7269: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5875Output_7270: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1395Output_7271: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5876Output_7272: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1396Output_7273: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5877Output_7274: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5879weight : std_logic_vector ( 22 downto 0 ) := "00111111001100010101001";

Signal ProductNode_POSIT5879Output_7276: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5881weight : std_logic_vector ( 22 downto 0 ) := "00111100110010101000000";

Signal ProductNode_POSIT5881Output_7278: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5882weight : std_logic_vector ( 22 downto 0 ) := "00111111111111001101010";

Signal ProductNode_POSIT5882Output_7279: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1397Output_7280: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5883Output_7281: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5888Output_7287: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5889weight : std_logic_vector ( 22 downto 0 ) := "00111100000000011010000";

Signal ProductNode_POSIT5889Output_7288: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5890weight : std_logic_vector ( 22 downto 0 ) := "00111111111111101111110";

Signal ProductNode_POSIT5890Output_7289: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1399Output_7290: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5891Output_7291: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5896Output_7297: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1401Output_7298: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5897Output_7299: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5906Output_7310: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5914Output_7320: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1406Output_7321: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5915Output_7322: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1407Output_7323: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5916Output_7324: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5948Output_7362: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5980Output_7400: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1420Output_7401: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5981Output_7402: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5983weight : std_logic_vector ( 22 downto 0 ) := "00111110100010010000110";

Signal ProductNode_POSIT5983Output_7404: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT5992Output_7415: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6000Output_7425: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1425Output_7426: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6001Output_7427: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6010Output_7438: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6018Output_7448: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1430Output_7449: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6019Output_7450: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1431Output_7451: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6020Output_7452: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6052Output_7490: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6084Output_7528: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1444Output_7529: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6085Output_7530: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1445Output_7531: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6086Output_7532: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6088weight : std_logic_vector ( 22 downto 0 ) := "00111111101001110101011";

Signal ProductNode_POSIT6088Output_7534: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6125Output_7582: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6157Output_7620: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6189Output_7658: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1469Output_7659: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6190Output_7660: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6192weight : std_logic_vector ( 22 downto 0 ) := "00111111110111011011110";

Signal ProductNode_POSIT6192Output_7662: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6229Output_7710: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6261Output_7748: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6293Output_7786: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1493Output_7787: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6294Output_7788: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1494Output_7789: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6295Output_7790: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1495Output_7791: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6296Output_7792: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6316Output_7817: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6334Output_7840: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1506Output_7841: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6335Output_7842: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6367Output_7880: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6399Output_7918: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1519Output_7919: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6400Output_7920: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6420Output_7945: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6438Output_7968: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1530Output_7969: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6439Output_7970: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6471Output_8008: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6503Output_8046: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1543Output_8047: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6504Output_8048: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1544Output_8049: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6505Output_8050: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6544Output_8100: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6576Output_8138: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6608Output_8176: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1568Output_8177: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6609Output_8178: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6648Output_8228: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6680Output_8266: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6712Output_8304: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1592Output_8305: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6713Output_8306: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1593Output_8307: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6714Output_8308: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1594Output_8309: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6715Output_8310: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1595Output_8311: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6716Output_8312: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1596Output_8313: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6717Output_8314: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1597Output_8315: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6718Output_8316: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1598Output_8317: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6719Output_8318: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6720weight : std_logic_vector ( 22 downto 0 ) := "00111111100000011111100";

Signal ProductNode_POSIT6720Output_8319: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6722weight : std_logic_vector ( 22 downto 0 ) := "00111111111100010100000";

Signal ProductNode_POSIT6722Output_8321: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6728weight : std_logic_vector ( 22 downto 0 ) := "00111111101110111111001";

Signal ProductNode_POSIT6728Output_8328: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6730weight : std_logic_vector ( 22 downto 0 ) := "00111111000010000001101";

Signal ProductNode_POSIT6730Output_8330: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1600Output_8331: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6731Output_8332: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6736weight : std_logic_vector ( 22 downto 0 ) := "00111111101110111111001";

Signal ProductNode_POSIT6736Output_8338: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6738weight : std_logic_vector ( 22 downto 0 ) := "00111111000010000001101";

Signal ProductNode_POSIT6738Output_8340: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1602Output_8341: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6739Output_8342: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1603Output_8343: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6740Output_8344: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6746weight : std_logic_vector ( 22 downto 0 ) := "00111111001000011011010";

Signal ProductNode_POSIT6746Output_8351: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6748weight : std_logic_vector ( 22 downto 0 ) := "00111111101011110010010";

Signal ProductNode_POSIT6748Output_8353: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1605Output_8354: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6749Output_8355: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6754weight : std_logic_vector ( 22 downto 0 ) := "00111111001000011011010";

Signal ProductNode_POSIT6754Output_8361: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6756weight : std_logic_vector ( 22 downto 0 ) := "00111111101011110010010";

Signal ProductNode_POSIT6756Output_8363: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1607Output_8364: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6757Output_8365: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1608Output_8366: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6758Output_8367: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1609Output_8368: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6759Output_8369: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6760weight : std_logic_vector ( 22 downto 0 ) := "00111111001010110111011";

Signal ProductNode_POSIT6760Output_8370: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6781Output_8394: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6782weight : std_logic_vector ( 22 downto 0 ) := "00111111011001110010110";

Signal ProductNode_POSIT6782Output_8395: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6786weight : std_logic_vector ( 22 downto 0 ) := "00111111111111001010111";

Signal ProductNode_POSIT6786Output_8400: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6790weight : std_logic_vector ( 22 downto 0 ) := "00111100110101000101000";

Signal ProductNode_POSIT6790Output_8405: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1615Output_8406: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6791Output_8407: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6792weight : std_logic_vector ( 22 downto 0 ) := "00111111101010100100010";

Signal ProductNode_POSIT6792Output_8408: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6813Output_8432: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6814weight : std_logic_vector ( 22 downto 0 ) := "00111111001001001110101";

Signal ProductNode_POSIT6814Output_8433: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6818weight : std_logic_vector ( 22 downto 0 ) := "00111111111110011110101";

Signal ProductNode_POSIT6818Output_8438: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6822weight : std_logic_vector ( 22 downto 0 ) := "00111101010000101001111";

Signal ProductNode_POSIT6822Output_8443: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1621Output_8444: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6823Output_8445: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1622Output_8446: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6824Output_8447: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6826weight : std_logic_vector ( 22 downto 0 ) := "00111111101110101011011";

Signal ProductNode_POSIT6826Output_8449: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6832weight : std_logic_vector ( 22 downto 0 ) := "00111111000111011011001";

Signal ProductNode_POSIT6832Output_8456: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6834weight : std_logic_vector ( 22 downto 0 ) := "00111111101100010010011";

Signal ProductNode_POSIT6834Output_8458: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1624Output_8459: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6835Output_8460: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6840weight : std_logic_vector ( 22 downto 0 ) := "00111111000111011011001";

Signal ProductNode_POSIT6840Output_8466: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6842weight : std_logic_vector ( 22 downto 0 ) := "00111111101100010010011";

Signal ProductNode_POSIT6842Output_8468: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1626Output_8469: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6843Output_8470: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1627Output_8471: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6844Output_8472: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6850weight : std_logic_vector ( 22 downto 0 ) := "00111110100101011101001";

Signal ProductNode_POSIT6850Output_8479: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6852weight : std_logic_vector ( 22 downto 0 ) := "00111111110110101000101";

Signal ProductNode_POSIT6852Output_8481: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1629Output_8482: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6853Output_8483: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6858weight : std_logic_vector ( 22 downto 0 ) := "00111110100101011101001";

Signal ProductNode_POSIT6858Output_8489: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6860weight : std_logic_vector ( 22 downto 0 ) := "00111111110110101000101";

Signal ProductNode_POSIT6860Output_8491: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1631Output_8492: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6861Output_8493: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1632Output_8494: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6862Output_8495: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1633Output_8496: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6863Output_8497: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6886weight : std_logic_vector ( 22 downto 0 ) := "00111111100011000110100";

Signal ProductNode_POSIT6886Output_8523: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6890weight : std_logic_vector ( 22 downto 0 ) := "00111111111110001110101";

Signal ProductNode_POSIT6890Output_8528: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6894weight : std_logic_vector ( 22 downto 0 ) := "00111101011000101001001";

Signal ProductNode_POSIT6894Output_8533: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1639Output_8534: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6895Output_8535: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6918weight : std_logic_vector ( 22 downto 0 ) := "00111111101011011000101";

Signal ProductNode_POSIT6918Output_8561: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6922weight : std_logic_vector ( 22 downto 0 ) := "00111111111111111110100";

Signal ProductNode_POSIT6922Output_8566: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6926weight : std_logic_vector ( 22 downto 0 ) := "00111010001101011110110";

Signal ProductNode_POSIT6926Output_8571: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1645Output_8572: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6927Output_8573: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1646Output_8574: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6928Output_8575: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1647Output_8576: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6929Output_8577: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6931weight : std_logic_vector ( 22 downto 0 ) := "00111101111010111110100";

Signal ProductNode_POSIT6931Output_8579: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6968Output_8627: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6995weight : std_logic_vector ( 22 downto 0 ) := "00111111110111110010101";

Signal ProductNode_POSIT6995Output_8658: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT6999weight : std_logic_vector ( 22 downto 0 ) := "00111110100000110101011";

Signal ProductNode_POSIT6999Output_8663: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1664Output_8664: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7000Output_8665: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7027weight : std_logic_vector ( 22 downto 0 ) := "00111111110010111011101";

Signal ProductNode_POSIT7027Output_8696: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7031weight : std_logic_vector ( 22 downto 0 ) := "00111110110100010001001";

Signal ProductNode_POSIT7031Output_8701: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1670Output_8702: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7032Output_8703: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1671Output_8704: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7033Output_8705: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7035weight : std_logic_vector ( 22 downto 0 ) := "00111111000010101001001";

Signal ProductNode_POSIT7035Output_8707: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7072Output_8755: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7099weight : std_logic_vector ( 22 downto 0 ) := "00111111101011011100110";

Signal ProductNode_POSIT7099Output_8786: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7103weight : std_logic_vector ( 22 downto 0 ) := "00111111001001000110010";

Signal ProductNode_POSIT7103Output_8791: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1688Output_8792: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7104Output_8793: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7131weight : std_logic_vector ( 22 downto 0 ) := "00111111011110011001000";

Signal ProductNode_POSIT7131Output_8824: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7135weight : std_logic_vector ( 22 downto 0 ) := "00111111100000110011011";

Signal ProductNode_POSIT7135Output_8829: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1694Output_8830: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7136Output_8831: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1695Output_8832: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7137Output_8833: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1696Output_8834: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7138Output_8835: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1697Output_8836: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7139Output_8837: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7159Output_8862: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7177Output_8885: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1708Output_8886: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7178Output_8887: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7200Output_8912: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7201weight : std_logic_vector ( 22 downto 0 ) := "00111110110100100010011";

Signal ProductNode_POSIT7201Output_8913: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7205weight : std_logic_vector ( 22 downto 0 ) := "00111111111011111111100";

Signal ProductNode_POSIT7205Output_8918: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7209weight : std_logic_vector ( 22 downto 0 ) := "00111110000000000011111";

Signal ProductNode_POSIT7209Output_8923: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1714Output_8924: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7210Output_8925: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7232Output_8950: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7233weight : std_logic_vector ( 22 downto 0 ) := "00111110001000001101101";

Signal ProductNode_POSIT7233Output_8951: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7237weight : std_logic_vector ( 22 downto 0 ) := "00111111111100000111010";

Signal ProductNode_POSIT7237Output_8956: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7241weight : std_logic_vector ( 22 downto 0 ) := "00111101111110001010101";

Signal ProductNode_POSIT7241Output_8961: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1720Output_8962: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7242Output_8963: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1721Output_8964: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7243Output_8965: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7263Output_8990: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7281Output_9013: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1732Output_9014: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7282Output_9015: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7305weight : std_logic_vector ( 22 downto 0 ) := "00111111110010110111011";

Signal ProductNode_POSIT7305Output_9041: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7309weight : std_logic_vector ( 22 downto 0 ) := "00111111111010111011111";

Signal ProductNode_POSIT7309Output_9046: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7313weight : std_logic_vector ( 22 downto 0 ) := "00111110001000100000100";

Signal ProductNode_POSIT7313Output_9051: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1738Output_9052: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7314Output_9053: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7337weight : std_logic_vector ( 22 downto 0 ) := "00111111111010111110010";

Signal ProductNode_POSIT7337Output_9079: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7341weight : std_logic_vector ( 22 downto 0 ) := "00111111111001110101001";

Signal ProductNode_POSIT7341Output_9084: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7345weight : std_logic_vector ( 22 downto 0 ) := "00111110010001010110100";

Signal ProductNode_POSIT7345Output_9089: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1744Output_9090: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7346Output_9091: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1745Output_9092: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7347Output_9093: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1746Output_9094: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7348Output_9095: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7387Output_9145: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7414weight : std_logic_vector ( 22 downto 0 ) := "00111111110000010101100";

Signal ProductNode_POSIT7414Output_9176: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7418weight : std_logic_vector ( 22 downto 0 ) := "00111110111110101001100";

Signal ProductNode_POSIT7418Output_9181: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1763Output_9182: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7419Output_9183: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7446weight : std_logic_vector ( 22 downto 0 ) := "00111111101111001010111";

Signal ProductNode_POSIT7446Output_9214: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7450weight : std_logic_vector ( 22 downto 0 ) := "00111111000001101010001";

Signal ProductNode_POSIT7450Output_9219: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1769Output_9220: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7451Output_9221: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1770Output_9222: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7452Output_9223: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7491Output_9273: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7518weight : std_logic_vector ( 22 downto 0 ) := "00111111100000110100110";

Signal ProductNode_POSIT7518Output_9304: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7522weight : std_logic_vector ( 22 downto 0 ) := "00111111011110010110011";

Signal ProductNode_POSIT7522Output_9309: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1787Output_9310: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7523Output_9311: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7550weight : std_logic_vector ( 22 downto 0 ) := "00111110111111110100001";

Signal ProductNode_POSIT7550Output_9342: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7554weight : std_logic_vector ( 22 downto 0 ) := "00111111110000000010111";

Signal ProductNode_POSIT7554Output_9347: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1793Output_9348: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7555Output_9349: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1794Output_9350: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7556Output_9351: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1795Output_9352: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7557Output_9353: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1796Output_9354: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7558Output_9355: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1797Output_9356: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7559Output_9357: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7561weight : std_logic_vector ( 22 downto 0 ) := "00111111111100010100000";

Signal ProductNode_POSIT7561Output_9359: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7570Output_9370: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7578Output_9380: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1802Output_9381: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7579Output_9382: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7588Output_9393: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7596Output_9403: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1807Output_9404: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7597Output_9405: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1808Output_9406: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7598Output_9407: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7620Output_9432: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7621weight : std_logic_vector ( 22 downto 0 ) := "00111111011001110010110";

Signal ProductNode_POSIT7621Output_9433: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7625weight : std_logic_vector ( 22 downto 0 ) := "00111111111111001010111";

Signal ProductNode_POSIT7625Output_9438: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7629weight : std_logic_vector ( 22 downto 0 ) := "00111100110101000101000";

Signal ProductNode_POSIT7629Output_9443: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1814Output_9444: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7630Output_9445: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7652Output_9470: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7653weight : std_logic_vector ( 22 downto 0 ) := "00111111001001001110101";

Signal ProductNode_POSIT7653Output_9471: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7657weight : std_logic_vector ( 22 downto 0 ) := "00111111111110011110101";

Signal ProductNode_POSIT7657Output_9476: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7661weight : std_logic_vector ( 22 downto 0 ) := "00111101010000101001111";

Signal ProductNode_POSIT7661Output_9481: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1820Output_9482: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7662Output_9483: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1821Output_9484: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7663Output_9485: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7665weight : std_logic_vector ( 22 downto 0 ) := "00111111101110101011011";

Signal ProductNode_POSIT7665Output_9487: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7674Output_9498: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7682Output_9508: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1826Output_9509: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7683Output_9510: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7692Output_9521: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7700Output_9531: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1831Output_9532: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7701Output_9533: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1832Output_9534: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7702Output_9535: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7725weight : std_logic_vector ( 22 downto 0 ) := "00111111100011000110100";

Signal ProductNode_POSIT7725Output_9561: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7729weight : std_logic_vector ( 22 downto 0 ) := "00111111111110001110101";

Signal ProductNode_POSIT7729Output_9566: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7733weight : std_logic_vector ( 22 downto 0 ) := "00111101011000101001001";

Signal ProductNode_POSIT7733Output_9571: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1838Output_9572: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7734Output_9573: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7757weight : std_logic_vector ( 22 downto 0 ) := "00111111101011011000101";

Signal ProductNode_POSIT7757Output_9599: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7761weight : std_logic_vector ( 22 downto 0 ) := "00111111111111111110100";

Signal ProductNode_POSIT7761Output_9604: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7765weight : std_logic_vector ( 22 downto 0 ) := "00111010001101011110110";

Signal ProductNode_POSIT7765Output_9609: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1844Output_9610: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7766Output_9611: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1845Output_9612: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7767Output_9613: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1846Output_9614: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7768Output_9615: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7770weight : std_logic_vector ( 22 downto 0 ) := "00111101111010111110100";

Signal ProductNode_POSIT7770Output_9617: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7807Output_9665: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7834weight : std_logic_vector ( 22 downto 0 ) := "00111111110111110010101";

Signal ProductNode_POSIT7834Output_9696: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7838weight : std_logic_vector ( 22 downto 0 ) := "00111110100000110101011";

Signal ProductNode_POSIT7838Output_9701: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1863Output_9702: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7839Output_9703: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7866weight : std_logic_vector ( 22 downto 0 ) := "00111111110010111011101";

Signal ProductNode_POSIT7866Output_9734: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7870weight : std_logic_vector ( 22 downto 0 ) := "00111110110100010001001";

Signal ProductNode_POSIT7870Output_9739: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1869Output_9740: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7871Output_9741: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1870Output_9742: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7872Output_9743: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7874weight : std_logic_vector ( 22 downto 0 ) := "00111111000010101001001";

Signal ProductNode_POSIT7874Output_9745: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7911Output_9793: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7938weight : std_logic_vector ( 22 downto 0 ) := "00111111101011011100110";

Signal ProductNode_POSIT7938Output_9824: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7942weight : std_logic_vector ( 22 downto 0 ) := "00111111001001000110010";

Signal ProductNode_POSIT7942Output_9829: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1887Output_9830: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7943Output_9831: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7970weight : std_logic_vector ( 22 downto 0 ) := "00111111011110011001000";

Signal ProductNode_POSIT7970Output_9862: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7974weight : std_logic_vector ( 22 downto 0 ) := "00111111100000110011011";

Signal ProductNode_POSIT7974Output_9867: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1893Output_9868: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7975Output_9869: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1894Output_9870: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7976Output_9871: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1895Output_9872: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7977Output_9873: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1896Output_9874: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7978Output_9875: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT7998Output_9900: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8016Output_9923: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1907Output_9924: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8017Output_9925: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8039Output_9950: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8040weight : std_logic_vector ( 22 downto 0 ) := "00111110110100100010011";

Signal ProductNode_POSIT8040Output_9951: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8044weight : std_logic_vector ( 22 downto 0 ) := "00111111111011111111100";

Signal ProductNode_POSIT8044Output_9956: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8048weight : std_logic_vector ( 22 downto 0 ) := "00111110000000000011111";

Signal ProductNode_POSIT8048Output_9961: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1913Output_9962: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8049Output_9963: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8071Output_9988: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8072weight : std_logic_vector ( 22 downto 0 ) := "00111110001000001101101";

Signal ProductNode_POSIT8072Output_9989: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8076weight : std_logic_vector ( 22 downto 0 ) := "00111111111100000111010";

Signal ProductNode_POSIT8076Output_9994: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8080weight : std_logic_vector ( 22 downto 0 ) := "00111101111110001010101";

Signal ProductNode_POSIT8080Output_9999: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1919Output_10000: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8081Output_10001: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1920Output_10002: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8082Output_10003: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8102Output_10028: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8120Output_10051: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1931Output_10052: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8121Output_10053: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8144weight : std_logic_vector ( 22 downto 0 ) := "00111111110010110111011";

Signal ProductNode_POSIT8144Output_10079: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8148weight : std_logic_vector ( 22 downto 0 ) := "00111111111010111011111";

Signal ProductNode_POSIT8148Output_10084: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8152weight : std_logic_vector ( 22 downto 0 ) := "00111110001000100000100";

Signal ProductNode_POSIT8152Output_10089: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1937Output_10090: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8153Output_10091: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8176weight : std_logic_vector ( 22 downto 0 ) := "00111111111010111110010";

Signal ProductNode_POSIT8176Output_10117: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8180weight : std_logic_vector ( 22 downto 0 ) := "00111111111001110101001";

Signal ProductNode_POSIT8180Output_10122: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8184weight : std_logic_vector ( 22 downto 0 ) := "00111110010001010110100";

Signal ProductNode_POSIT8184Output_10127: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1943Output_10128: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8185Output_10129: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1944Output_10130: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8186Output_10131: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1945Output_10132: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8187Output_10133: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8226Output_10183: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8253weight : std_logic_vector ( 22 downto 0 ) := "00111111110000010101100";

Signal ProductNode_POSIT8253Output_10214: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8257weight : std_logic_vector ( 22 downto 0 ) := "00111110111110101001100";

Signal ProductNode_POSIT8257Output_10219: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1962Output_10220: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8258Output_10221: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8285weight : std_logic_vector ( 22 downto 0 ) := "00111111101111001010111";

Signal ProductNode_POSIT8285Output_10252: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8289weight : std_logic_vector ( 22 downto 0 ) := "00111111000001101010001";

Signal ProductNode_POSIT8289Output_10257: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1968Output_10258: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8290Output_10259: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1969Output_10260: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8291Output_10261: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8330Output_10311: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8357weight : std_logic_vector ( 22 downto 0 ) := "00111111100000110100110";

Signal ProductNode_POSIT8357Output_10342: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8361weight : std_logic_vector ( 22 downto 0 ) := "00111111011110010110011";

Signal ProductNode_POSIT8361Output_10347: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1986Output_10348: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8362Output_10349: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8389weight : std_logic_vector ( 22 downto 0 ) := "00111110111111110100001";

Signal ProductNode_POSIT8389Output_10380: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8393weight : std_logic_vector ( 22 downto 0 ) := "00111111110000000010111";

Signal ProductNode_POSIT8393Output_10385: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1992Output_10386: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8394Output_10387: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1993Output_10388: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8395Output_10389: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1994Output_10390: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8396Output_10391: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1995Output_10392: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8397Output_10393: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1996Output_10394: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8398Output_10395: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1997Output_10396: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8399Output_10397: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8401weight : std_logic_vector ( 22 downto 0 ) := "00111111011001010011000";

Signal ProductNode_POSIT8401Output_10399: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8407weight : std_logic_vector ( 22 downto 0 ) := "00111111001111110111000";

Signal ProductNode_POSIT8407Output_10406: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8409weight : std_logic_vector ( 22 downto 0 ) := "00111111101000000100011";

Signal ProductNode_POSIT8409Output_10408: std_logic_vector (22 downto 0);
Signal SumNode_POSIT1999Output_10409: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8410Output_10410: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8415weight : std_logic_vector ( 22 downto 0 ) := "00111111001111110111000";

Signal ProductNode_POSIT8415Output_10416: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8417weight : std_logic_vector ( 22 downto 0 ) := "00111111101000000100011";

Signal ProductNode_POSIT8417Output_10418: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2001Output_10419: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8418Output_10420: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2002Output_10421: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8419Output_10422: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8425weight : std_logic_vector ( 22 downto 0 ) := "00111110100100101101001";

Signal ProductNode_POSIT8425Output_10429: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8427weight : std_logic_vector ( 22 downto 0 ) := "00111111110110110100101";

Signal ProductNode_POSIT8427Output_10431: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2004Output_10432: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8428Output_10433: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8433weight : std_logic_vector ( 22 downto 0 ) := "00111110100100101101001";

Signal ProductNode_POSIT8433Output_10439: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8435weight : std_logic_vector ( 22 downto 0 ) := "00111111110110110100101";

Signal ProductNode_POSIT8435Output_10441: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2006Output_10442: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8436Output_10443: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2007Output_10444: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8437Output_10445: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2008Output_10446: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8438Output_10447: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8465weight : std_logic_vector ( 22 downto 0 ) := "00111111111111001010111";

Signal ProductNode_POSIT8465Output_10478: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8469weight : std_logic_vector ( 22 downto 0 ) := "00111100110101000101000";

Signal ProductNode_POSIT8469Output_10483: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2014Output_10484: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8470Output_10485: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8497weight : std_logic_vector ( 22 downto 0 ) := "00111111111110011110101";

Signal ProductNode_POSIT8497Output_10516: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8501weight : std_logic_vector ( 22 downto 0 ) := "00111101010000101001111";

Signal ProductNode_POSIT8501Output_10521: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2020Output_10522: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8502Output_10523: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2021Output_10524: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8503Output_10525: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8505weight : std_logic_vector ( 22 downto 0 ) := "00111110100010000010110";

Signal ProductNode_POSIT8505Output_10527: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8511weight : std_logic_vector ( 22 downto 0 ) := "00111110101001001010011";

Signal ProductNode_POSIT8511Output_10534: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8513weight : std_logic_vector ( 22 downto 0 ) := "00111111110101101101011";

Signal ProductNode_POSIT8513Output_10536: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2023Output_10537: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8514Output_10538: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8519weight : std_logic_vector ( 22 downto 0 ) := "00111110101001001010011";

Signal ProductNode_POSIT8519Output_10544: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8521weight : std_logic_vector ( 22 downto 0 ) := "00111111110101101101011";

Signal ProductNode_POSIT8521Output_10546: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2025Output_10547: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8522Output_10548: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2026Output_10549: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8523Output_10550: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8529weight : std_logic_vector ( 22 downto 0 ) := "00111101000101011011011";

Signal ProductNode_POSIT8529Output_10557: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8531weight : std_logic_vector ( 22 downto 0 ) := "00111111111110110101001";

Signal ProductNode_POSIT8531Output_10559: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2028Output_10560: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8532Output_10561: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8537weight : std_logic_vector ( 22 downto 0 ) := "00111101000101011011011";

Signal ProductNode_POSIT8537Output_10567: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8539weight : std_logic_vector ( 22 downto 0 ) := "00111111111110110101001";

Signal ProductNode_POSIT8539Output_10569: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2030Output_10570: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8540Output_10571: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2031Output_10572: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8541Output_10573: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2032Output_10574: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8542Output_10575: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8569weight : std_logic_vector ( 22 downto 0 ) := "00111111111110001110101";

Signal ProductNode_POSIT8569Output_10606: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8573weight : std_logic_vector ( 22 downto 0 ) := "00111101011000101001001";

Signal ProductNode_POSIT8573Output_10611: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2038Output_10612: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8574Output_10613: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8601weight : std_logic_vector ( 22 downto 0 ) := "00111111111111111110100";

Signal ProductNode_POSIT8601Output_10644: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8605weight : std_logic_vector ( 22 downto 0 ) := "00111010001101011110110";

Signal ProductNode_POSIT8605Output_10649: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2044Output_10650: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8606Output_10651: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2045Output_10652: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8607Output_10653: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2046Output_10654: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8608Output_10655: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8610weight : std_logic_vector ( 22 downto 0 ) := "00111111100011010110011";

Signal ProductNode_POSIT8610Output_10657: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8647Output_10705: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8674weight : std_logic_vector ( 22 downto 0 ) := "00111111110111110010101";

Signal ProductNode_POSIT8674Output_10736: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8678weight : std_logic_vector ( 22 downto 0 ) := "00111110100000110101011";

Signal ProductNode_POSIT8678Output_10741: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2063Output_10742: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8679Output_10743: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8706weight : std_logic_vector ( 22 downto 0 ) := "00111111110010111011101";

Signal ProductNode_POSIT8706Output_10774: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8710weight : std_logic_vector ( 22 downto 0 ) := "00111110110100010001001";

Signal ProductNode_POSIT8710Output_10779: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2069Output_10780: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8711Output_10781: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2070Output_10782: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8712Output_10783: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8714weight : std_logic_vector ( 22 downto 0 ) := "00111111110111011111010";

Signal ProductNode_POSIT8714Output_10785: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8751Output_10833: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8778weight : std_logic_vector ( 22 downto 0 ) := "00111111101011011100110";

Signal ProductNode_POSIT8778Output_10864: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8782weight : std_logic_vector ( 22 downto 0 ) := "00111111001001000110010";

Signal ProductNode_POSIT8782Output_10869: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2087Output_10870: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8783Output_10871: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8810weight : std_logic_vector ( 22 downto 0 ) := "00111111011110011001000";

Signal ProductNode_POSIT8810Output_10902: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8814weight : std_logic_vector ( 22 downto 0 ) := "00111111100000110011011";

Signal ProductNode_POSIT8814Output_10907: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2093Output_10908: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8815Output_10909: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2094Output_10910: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8816Output_10911: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2095Output_10912: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8817Output_10913: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2096Output_10914: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8818Output_10915: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8838Output_10940: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8856Output_10963: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2107Output_10964: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8857Output_10965: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8884weight : std_logic_vector ( 22 downto 0 ) := "00111111111011111111100";

Signal ProductNode_POSIT8884Output_10996: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8888weight : std_logic_vector ( 22 downto 0 ) := "00111110000000000011111";

Signal ProductNode_POSIT8888Output_11001: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2113Output_11002: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8889Output_11003: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8916weight : std_logic_vector ( 22 downto 0 ) := "00111111111100000111010";

Signal ProductNode_POSIT8916Output_11034: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8920weight : std_logic_vector ( 22 downto 0 ) := "00111101111110001010101";

Signal ProductNode_POSIT8920Output_11039: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2119Output_11040: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8921Output_11041: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2120Output_11042: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8922Output_11043: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8942Output_11068: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8960Output_11091: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2131Output_11092: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8961Output_11093: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8988weight : std_logic_vector ( 22 downto 0 ) := "00111111111010111011111";

Signal ProductNode_POSIT8988Output_11124: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8992weight : std_logic_vector ( 22 downto 0 ) := "00111110001000100000100";

Signal ProductNode_POSIT8992Output_11129: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2137Output_11130: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT8993Output_11131: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9020weight : std_logic_vector ( 22 downto 0 ) := "00111111111001110101001";

Signal ProductNode_POSIT9020Output_11162: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9024weight : std_logic_vector ( 22 downto 0 ) := "00111110010001010110100";

Signal ProductNode_POSIT9024Output_11167: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2143Output_11168: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9025Output_11169: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2144Output_11170: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9026Output_11171: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2145Output_11172: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9027Output_11173: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9066Output_11223: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9093weight : std_logic_vector ( 22 downto 0 ) := "00111111110000010101100";

Signal ProductNode_POSIT9093Output_11254: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9097weight : std_logic_vector ( 22 downto 0 ) := "00111110111110101001100";

Signal ProductNode_POSIT9097Output_11259: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2162Output_11260: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9098Output_11261: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9125weight : std_logic_vector ( 22 downto 0 ) := "00111111101111001010111";

Signal ProductNode_POSIT9125Output_11292: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9129weight : std_logic_vector ( 22 downto 0 ) := "00111111000001101010001";

Signal ProductNode_POSIT9129Output_11297: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2168Output_11298: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9130Output_11299: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2169Output_11300: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9131Output_11301: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9170Output_11351: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9197weight : std_logic_vector ( 22 downto 0 ) := "00111111100000110100110";

Signal ProductNode_POSIT9197Output_11382: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9201weight : std_logic_vector ( 22 downto 0 ) := "00111111011110010110011";

Signal ProductNode_POSIT9201Output_11387: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2186Output_11388: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9202Output_11389: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9229weight : std_logic_vector ( 22 downto 0 ) := "00111110111111110100001";

Signal ProductNode_POSIT9229Output_11420: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9233weight : std_logic_vector ( 22 downto 0 ) := "00111111110000000010111";

Signal ProductNode_POSIT9233Output_11425: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2192Output_11426: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9234Output_11427: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2193Output_11428: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9235Output_11429: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2194Output_11430: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9236Output_11431: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2195Output_11432: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9237Output_11433: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2196Output_11434: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9238Output_11435: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9240weight : std_logic_vector ( 22 downto 0 ) := "00111111011001010011000";

Signal ProductNode_POSIT9240Output_11437: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9249Output_11448: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9257Output_11458: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2201Output_11459: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9258Output_11460: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9267Output_11471: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9275Output_11481: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2206Output_11482: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9276Output_11483: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2207Output_11484: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9277Output_11485: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9304weight : std_logic_vector ( 22 downto 0 ) := "00111111111111001010111";

Signal ProductNode_POSIT9304Output_11516: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9308weight : std_logic_vector ( 22 downto 0 ) := "00111100110101000101000";

Signal ProductNode_POSIT9308Output_11521: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2213Output_11522: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9309Output_11523: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9336weight : std_logic_vector ( 22 downto 0 ) := "00111111111110011110101";

Signal ProductNode_POSIT9336Output_11554: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9340weight : std_logic_vector ( 22 downto 0 ) := "00111101010000101001111";

Signal ProductNode_POSIT9340Output_11559: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2219Output_11560: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9341Output_11561: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2220Output_11562: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9342Output_11563: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9344weight : std_logic_vector ( 22 downto 0 ) := "00111110100010000010110";

Signal ProductNode_POSIT9344Output_11565: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9353Output_11576: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9361Output_11586: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2225Output_11587: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9362Output_11588: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9371Output_11599: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9379Output_11609: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2230Output_11610: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9380Output_11611: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2231Output_11612: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9381Output_11613: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9408weight : std_logic_vector ( 22 downto 0 ) := "00111111111110001110101";

Signal ProductNode_POSIT9408Output_11644: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9412weight : std_logic_vector ( 22 downto 0 ) := "00111101011000101001001";

Signal ProductNode_POSIT9412Output_11649: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2237Output_11650: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9413Output_11651: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9440weight : std_logic_vector ( 22 downto 0 ) := "00111111111111111110100";

Signal ProductNode_POSIT9440Output_11682: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9444weight : std_logic_vector ( 22 downto 0 ) := "00111010001101011110110";

Signal ProductNode_POSIT9444Output_11687: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2243Output_11688: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9445Output_11689: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2244Output_11690: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9446Output_11691: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2245Output_11692: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9447Output_11693: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9449weight : std_logic_vector ( 22 downto 0 ) := "00111111100011010110011";

Signal ProductNode_POSIT9449Output_11695: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9486Output_11743: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9513weight : std_logic_vector ( 22 downto 0 ) := "00111111110111110010101";

Signal ProductNode_POSIT9513Output_11774: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9517weight : std_logic_vector ( 22 downto 0 ) := "00111110100000110101011";

Signal ProductNode_POSIT9517Output_11779: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2262Output_11780: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9518Output_11781: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9545weight : std_logic_vector ( 22 downto 0 ) := "00111111110010111011101";

Signal ProductNode_POSIT9545Output_11812: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9549weight : std_logic_vector ( 22 downto 0 ) := "00111110110100010001001";

Signal ProductNode_POSIT9549Output_11817: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2268Output_11818: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9550Output_11819: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2269Output_11820: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9551Output_11821: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9553weight : std_logic_vector ( 22 downto 0 ) := "00111111110111011111010";

Signal ProductNode_POSIT9553Output_11823: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9590Output_11871: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9617weight : std_logic_vector ( 22 downto 0 ) := "00111111101011011100110";

Signal ProductNode_POSIT9617Output_11902: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9621weight : std_logic_vector ( 22 downto 0 ) := "00111111001001000110010";

Signal ProductNode_POSIT9621Output_11907: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2286Output_11908: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9622Output_11909: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9649weight : std_logic_vector ( 22 downto 0 ) := "00111111011110011001000";

Signal ProductNode_POSIT9649Output_11940: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9653weight : std_logic_vector ( 22 downto 0 ) := "00111111100000110011011";

Signal ProductNode_POSIT9653Output_11945: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2292Output_11946: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9654Output_11947: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2293Output_11948: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9655Output_11949: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2294Output_11950: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9656Output_11951: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2295Output_11952: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9657Output_11953: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9677Output_11978: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9695Output_12001: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2306Output_12002: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9696Output_12003: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9723weight : std_logic_vector ( 22 downto 0 ) := "00111111111011111111100";

Signal ProductNode_POSIT9723Output_12034: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9727weight : std_logic_vector ( 22 downto 0 ) := "00111110000000000011111";

Signal ProductNode_POSIT9727Output_12039: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2312Output_12040: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9728Output_12041: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9755weight : std_logic_vector ( 22 downto 0 ) := "00111111111100000111010";

Signal ProductNode_POSIT9755Output_12072: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9759weight : std_logic_vector ( 22 downto 0 ) := "00111101111110001010101";

Signal ProductNode_POSIT9759Output_12077: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2318Output_12078: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9760Output_12079: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2319Output_12080: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9761Output_12081: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9781Output_12106: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9799Output_12129: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2330Output_12130: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9800Output_12131: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9827weight : std_logic_vector ( 22 downto 0 ) := "00111111111010111011111";

Signal ProductNode_POSIT9827Output_12162: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9831weight : std_logic_vector ( 22 downto 0 ) := "00111110001000100000100";

Signal ProductNode_POSIT9831Output_12167: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2336Output_12168: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9832Output_12169: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9859weight : std_logic_vector ( 22 downto 0 ) := "00111111111001110101001";

Signal ProductNode_POSIT9859Output_12200: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9863weight : std_logic_vector ( 22 downto 0 ) := "00111110010001010110100";

Signal ProductNode_POSIT9863Output_12205: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2342Output_12206: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9864Output_12207: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2343Output_12208: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9865Output_12209: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2344Output_12210: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9866Output_12211: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9905Output_12261: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9932weight : std_logic_vector ( 22 downto 0 ) := "00111111110000010101100";

Signal ProductNode_POSIT9932Output_12292: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9936weight : std_logic_vector ( 22 downto 0 ) := "00111110111110101001100";

Signal ProductNode_POSIT9936Output_12297: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2361Output_12298: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9937Output_12299: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9964weight : std_logic_vector ( 22 downto 0 ) := "00111111101111001010111";

Signal ProductNode_POSIT9964Output_12330: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9968weight : std_logic_vector ( 22 downto 0 ) := "00111111000001101010001";

Signal ProductNode_POSIT9968Output_12335: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2367Output_12336: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9969Output_12337: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2368Output_12338: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT9970Output_12339: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10009Output_12389: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10036weight : std_logic_vector ( 22 downto 0 ) := "00111111100000110100110";

Signal ProductNode_POSIT10036Output_12420: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10040weight : std_logic_vector ( 22 downto 0 ) := "00111111011110010110011";

Signal ProductNode_POSIT10040Output_12425: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2385Output_12426: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10041Output_12427: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10068weight : std_logic_vector ( 22 downto 0 ) := "00111110111111110100001";

Signal ProductNode_POSIT10068Output_12458: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10072weight : std_logic_vector ( 22 downto 0 ) := "00111111110000000010111";

Signal ProductNode_POSIT10072Output_12463: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2391Output_12464: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10073Output_12465: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2392Output_12466: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10074Output_12467: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2393Output_12468: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10075Output_12469: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2394Output_12470: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10076Output_12471: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2395Output_12472: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10077Output_12473: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2396Output_12474: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10078Output_12475: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2397Output_12476: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10079Output_12477: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10081weight : std_logic_vector ( 22 downto 0 ) := "00111111110100010010001";

Signal ProductNode_POSIT10081Output_12479: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10090Output_12490: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10098Output_12500: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2402Output_12501: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10099Output_12502: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10108Output_12513: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10116Output_12523: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2407Output_12524: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10117Output_12525: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2408Output_12526: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10118Output_12527: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10140Output_12552: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10141weight : std_logic_vector ( 22 downto 0 ) := "00111111011001110010110";

Signal ProductNode_POSIT10141Output_12553: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10150Output_12565: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10172Output_12590: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10173weight : std_logic_vector ( 22 downto 0 ) := "00111111001001001110101";

Signal ProductNode_POSIT10173Output_12591: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10182Output_12603: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2421Output_12604: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10183Output_12605: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10185weight : std_logic_vector ( 22 downto 0 ) := "00111111100011001010011";

Signal ProductNode_POSIT10185Output_12607: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10194Output_12618: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10202Output_12628: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2426Output_12629: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10203Output_12630: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10212Output_12641: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10220Output_12651: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2431Output_12652: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10221Output_12653: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2432Output_12654: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10222Output_12655: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10245weight : std_logic_vector ( 22 downto 0 ) := "00111111100011000110100";

Signal ProductNode_POSIT10245Output_12681: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10254Output_12693: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10277weight : std_logic_vector ( 22 downto 0 ) := "00111111101011011000101";

Signal ProductNode_POSIT10277Output_12719: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10286Output_12731: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2445Output_12732: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10287Output_12733: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2446Output_12734: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10288Output_12735: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10290weight : std_logic_vector ( 22 downto 0 ) := "00111110101110110111010";

Signal ProductNode_POSIT10290Output_12737: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10327Output_12785: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10359Output_12823: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10391Output_12861: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2470Output_12862: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10392Output_12863: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10394weight : std_logic_vector ( 22 downto 0 ) := "00111111011001101011001";

Signal ProductNode_POSIT10394Output_12865: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10431Output_12913: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10463Output_12951: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10495Output_12989: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2494Output_12990: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10496Output_12991: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2495Output_12992: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10497Output_12993: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2496Output_12994: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10498Output_12995: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10518Output_13020: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10536Output_13043: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2507Output_13044: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10537Output_13045: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10559Output_13070: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10560weight : std_logic_vector ( 22 downto 0 ) := "00111110110100100010011";

Signal ProductNode_POSIT10560Output_13071: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10569Output_13083: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10591Output_13108: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10592weight : std_logic_vector ( 22 downto 0 ) := "00111110001000001101101";

Signal ProductNode_POSIT10592Output_13109: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10601Output_13121: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2520Output_13122: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10602Output_13123: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10622Output_13148: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10640Output_13171: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2531Output_13172: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10641Output_13173: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10664weight : std_logic_vector ( 22 downto 0 ) := "00111111110010110111011";

Signal ProductNode_POSIT10664Output_13199: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10673Output_13211: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10696weight : std_logic_vector ( 22 downto 0 ) := "00111111111010111110010";

Signal ProductNode_POSIT10696Output_13237: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10705Output_13249: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2544Output_13250: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10706Output_13251: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2545Output_13252: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10707Output_13253: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10746Output_13303: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10778Output_13341: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10810Output_13379: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2569Output_13380: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10811Output_13381: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10850Output_13431: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10882Output_13469: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10914Output_13507: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2593Output_13508: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10915Output_13509: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2594Output_13510: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10916Output_13511: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2595Output_13512: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10917Output_13513: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2596Output_13514: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10918Output_13515: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10920weight : std_logic_vector ( 22 downto 0 ) := "00111111110100010010001";

Signal ProductNode_POSIT10920Output_13517: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10929Output_13528: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10937Output_13538: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2601Output_13539: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10938Output_13540: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10947Output_13551: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10955Output_13561: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2606Output_13562: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10956Output_13563: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2607Output_13564: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10957Output_13565: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10979Output_13590: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10980weight : std_logic_vector ( 22 downto 0 ) := "00111111011001110010110";

Signal ProductNode_POSIT10980Output_13591: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT10989Output_13603: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11011Output_13628: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11012weight : std_logic_vector ( 22 downto 0 ) := "00111111001001001110101";

Signal ProductNode_POSIT11012Output_13629: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11021Output_13641: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2620Output_13642: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11022Output_13643: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11024weight : std_logic_vector ( 22 downto 0 ) := "00111111100011001010011";

Signal ProductNode_POSIT11024Output_13645: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11033Output_13656: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11041Output_13666: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2625Output_13667: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11042Output_13668: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11051Output_13679: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11059Output_13689: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2630Output_13690: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11060Output_13691: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2631Output_13692: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11061Output_13693: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11084weight : std_logic_vector ( 22 downto 0 ) := "00111111100011000110100";

Signal ProductNode_POSIT11084Output_13719: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11093Output_13731: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11116weight : std_logic_vector ( 22 downto 0 ) := "00111111101011011000101";

Signal ProductNode_POSIT11116Output_13757: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11125Output_13769: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2644Output_13770: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11126Output_13771: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2645Output_13772: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11127Output_13773: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11129weight : std_logic_vector ( 22 downto 0 ) := "00111110101110110111010";

Signal ProductNode_POSIT11129Output_13775: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11166Output_13823: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11198Output_13861: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11230Output_13899: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2669Output_13900: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11231Output_13901: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11233weight : std_logic_vector ( 22 downto 0 ) := "00111111011001101011001";

Signal ProductNode_POSIT11233Output_13903: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11270Output_13951: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11302Output_13989: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11334Output_14027: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2693Output_14028: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11335Output_14029: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2694Output_14030: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11336Output_14031: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2695Output_14032: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11337Output_14033: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11357Output_14058: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11375Output_14081: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2706Output_14082: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11376Output_14083: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11398Output_14108: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11399weight : std_logic_vector ( 22 downto 0 ) := "00111110110100100010011";

Signal ProductNode_POSIT11399Output_14109: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11408Output_14121: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11430Output_14146: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11431weight : std_logic_vector ( 22 downto 0 ) := "00111110001000001101101";

Signal ProductNode_POSIT11431Output_14147: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11440Output_14159: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2719Output_14160: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11441Output_14161: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11461Output_14186: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11479Output_14209: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2730Output_14210: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11480Output_14211: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11503weight : std_logic_vector ( 22 downto 0 ) := "00111111110010110111011";

Signal ProductNode_POSIT11503Output_14237: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11512Output_14249: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11535weight : std_logic_vector ( 22 downto 0 ) := "00111111111010111110010";

Signal ProductNode_POSIT11535Output_14275: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11544Output_14287: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2743Output_14288: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11545Output_14289: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2744Output_14290: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11546Output_14291: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11585Output_14341: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11617Output_14379: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11649Output_14417: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2768Output_14418: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11650Output_14419: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11689Output_14469: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11721Output_14507: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11753Output_14545: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2792Output_14546: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11754Output_14547: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2793Output_14548: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11755Output_14549: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2794Output_14550: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11756Output_14551: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2795Output_14552: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11757Output_14553: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2796Output_14554: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11758Output_14555: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11760weight : std_logic_vector ( 22 downto 0 ) := "00111111000101001000010";

Signal ProductNode_POSIT11760Output_14557: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11769Output_14568: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11777Output_14578: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2801Output_14579: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11778Output_14580: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11787Output_14591: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11795Output_14601: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2806Output_14602: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11796Output_14603: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2807Output_14604: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11797Output_14605: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11829Output_14643: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11861Output_14681: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2820Output_14682: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11862Output_14683: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11864weight : std_logic_vector ( 22 downto 0 ) := "00111101100101010010010";

Signal ProductNode_POSIT11864Output_14685: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11873Output_14696: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11881Output_14706: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2825Output_14707: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11882Output_14708: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11891Output_14719: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11899Output_14729: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2830Output_14730: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11900Output_14731: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2831Output_14732: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11901Output_14733: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11933Output_14771: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11965Output_14809: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2844Output_14810: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11966Output_14811: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2845Output_14812: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11967Output_14813: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT11969weight : std_logic_vector ( 22 downto 0 ) := "00111111101101011011110";

Signal ProductNode_POSIT11969Output_14815: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT12006Output_14863: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT12038Output_14901: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT12070Output_14939: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2869Output_14940: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT12071Output_14941: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT12073weight : std_logic_vector ( 22 downto 0 ) := "00111111111101101010110";

Signal ProductNode_POSIT12073Output_14943: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT12110Output_14991: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT12142Output_15029: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT12174Output_15067: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2893Output_15068: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT12175Output_15069: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2894Output_15070: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT12176Output_15071: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2895Output_15072: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT12177Output_15073: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT12197Output_15098: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT12215Output_15121: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2906Output_15122: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT12216Output_15123: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT12248Output_15161: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT12280Output_15199: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2919Output_15200: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT12281Output_15201: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT12301Output_15226: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT12319Output_15249: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2930Output_15250: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT12320Output_15251: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT12352Output_15289: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT12384Output_15327: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2943Output_15328: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT12385Output_15329: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2944Output_15330: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT12386Output_15331: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT12425Output_15381: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT12457Output_15419: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT12489Output_15457: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2968Output_15458: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT12490Output_15459: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT12529Output_15509: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT12561Output_15547: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT12593Output_15585: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2992Output_15586: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT12594Output_15587: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2993Output_15588: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT12595Output_15589: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2994Output_15590: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT12596Output_15591: std_logic_vector (22 downto 0);
Signal SumNode_POSIT2995Output_15592: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT12597Output_15593: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT12599weight : std_logic_vector ( 22 downto 0 ) := "00111111000101001000010";

Signal ProductNode_POSIT12599Output_15595: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT12608Output_15606: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT12616Output_15616: std_logic_vector (22 downto 0);
Signal SumNode_POSIT3000Output_15617: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT12617Output_15618: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT12626Output_15629: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT12634Output_15639: std_logic_vector (22 downto 0);
Signal SumNode_POSIT3005Output_15640: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT12635Output_15641: std_logic_vector (22 downto 0);
Signal SumNode_POSIT3006Output_15642: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT12636Output_15643: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT12668Output_15681: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT12700Output_15719: std_logic_vector (22 downto 0);
Signal SumNode_POSIT3019Output_15720: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT12701Output_15721: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT12703weight : std_logic_vector ( 22 downto 0 ) := "00111101100101010010010";

Signal ProductNode_POSIT12703Output_15723: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT12712Output_15734: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT12720Output_15744: std_logic_vector (22 downto 0);
Signal SumNode_POSIT3024Output_15745: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT12721Output_15746: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT12730Output_15757: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT12738Output_15767: std_logic_vector (22 downto 0);
Signal SumNode_POSIT3029Output_15768: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT12739Output_15769: std_logic_vector (22 downto 0);
Signal SumNode_POSIT3030Output_15770: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT12740Output_15771: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT12772Output_15809: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT12804Output_15847: std_logic_vector (22 downto 0);
Signal SumNode_POSIT3043Output_15848: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT12805Output_15849: std_logic_vector (22 downto 0);
Signal SumNode_POSIT3044Output_15850: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT12806Output_15851: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT12808weight : std_logic_vector ( 22 downto 0 ) := "00111111101101011011110";

Signal ProductNode_POSIT12808Output_15853: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT12845Output_15901: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT12877Output_15939: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT12909Output_15977: std_logic_vector (22 downto 0);
Signal SumNode_POSIT3068Output_15978: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT12910Output_15979: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT12912weight : std_logic_vector ( 22 downto 0 ) := "00111111111101101010110";

Signal ProductNode_POSIT12912Output_15981: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT12949Output_16029: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT12981Output_16067: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT13013Output_16105: std_logic_vector (22 downto 0);
Signal SumNode_POSIT3092Output_16106: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT13014Output_16107: std_logic_vector (22 downto 0);
Signal SumNode_POSIT3093Output_16108: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT13015Output_16109: std_logic_vector (22 downto 0);
Signal SumNode_POSIT3094Output_16110: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT13016Output_16111: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT13036Output_16136: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT13054Output_16159: std_logic_vector (22 downto 0);
Signal SumNode_POSIT3105Output_16160: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT13055Output_16161: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT13087Output_16199: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT13119Output_16237: std_logic_vector (22 downto 0);
Signal SumNode_POSIT3118Output_16238: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT13120Output_16239: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT13140Output_16264: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT13158Output_16287: std_logic_vector (22 downto 0);
Signal SumNode_POSIT3129Output_16288: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT13159Output_16289: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT13191Output_16327: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT13223Output_16365: std_logic_vector (22 downto 0);
Signal SumNode_POSIT3142Output_16366: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT13224Output_16367: std_logic_vector (22 downto 0);
Signal SumNode_POSIT3143Output_16368: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT13225Output_16369: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT13264Output_16419: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT13296Output_16457: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT13328Output_16495: std_logic_vector (22 downto 0);
Signal SumNode_POSIT3167Output_16496: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT13329Output_16497: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT13368Output_16547: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT13400Output_16585: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT13432Output_16623: std_logic_vector (22 downto 0);
Signal SumNode_POSIT3191Output_16624: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT13433Output_16625: std_logic_vector (22 downto 0);
Signal SumNode_POSIT3192Output_16626: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT13434Output_16627: std_logic_vector (22 downto 0);
Signal SumNode_POSIT3193Output_16628: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT13435Output_16629: std_logic_vector (22 downto 0);
Signal SumNode_POSIT3194Output_16630: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT13436Output_16631: std_logic_vector (22 downto 0);
Signal SumNode_POSIT3195Output_16632: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT13437Output_16633: std_logic_vector (22 downto 0);
Signal SumNode_POSIT3196Output_16634: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT13438Output_16635: std_logic_vector (22 downto 0);
Signal SumNode_POSIT3197Output_16636: std_logic_vector (22 downto 0);
Signal ProductNode_POSIT13439Output_16637: std_logic_vector (22 downto 0);
Signal SumNode_POSIT3198Output_16638: std_logic_vector (22 downto 0);

 
begin 
ProductNode_POSIT0: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT0weight,v9,ProductNode_POSIT0Output_0);

ProductNode_POSIT1: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1weight,v11,ProductNode_POSIT1Output_1);

ProductNode_POSIT2: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT2weight,ProductNode_POSIT1Output_1,ProductNode_POSIT2Output_2);

ProductNode_POSIT3: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT3weight,v2,ProductNode_POSIT3Output_3);

ProductNode_POSIT4: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT4weight,v7,ProductNode_POSIT4Output_4);

ProductNode_POSIT5: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT5weight,vb7,ProductNode_POSIT5Output_5);

SumNode_POSIT0: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT5Output_5,ProductNode_POSIT4Output_4,SumNode_POSIT0Output_6);

ProductNode_POSIT6: entity work.PositMult_23_6_comb_uid2(arch)
port map(v1,SumNode_POSIT0Output_6,ProductNode_POSIT6Output_7);

ProductNode_POSIT7: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT7weight,v8,ProductNode_POSIT7Output_8);

ProductNode_POSIT8: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT8weight,ProductNode_POSIT7Output_8,ProductNode_POSIT8Output_9);

ProductNode_POSIT9: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT9weight,vb8,ProductNode_POSIT9Output_10);

ProductNode_POSIT10: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT10weight,ProductNode_POSIT9Output_10,ProductNode_POSIT10Output_11);

SumNode_POSIT1: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT10Output_11,ProductNode_POSIT8Output_9,SumNode_POSIT1Output_12);

ProductNode_POSIT11: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1Output_12,ProductNode_POSIT6Output_7,ProductNode_POSIT11Output_13);

ProductNode_POSIT12: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT12weight,v7,ProductNode_POSIT12Output_14);

ProductNode_POSIT13: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT13weight,vb7,ProductNode_POSIT13Output_15);

SumNode_POSIT2: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT13Output_15,ProductNode_POSIT12Output_14,SumNode_POSIT2Output_16);

ProductNode_POSIT14: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb1,SumNode_POSIT2Output_16,ProductNode_POSIT14Output_17);

ProductNode_POSIT15: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT15weight,v8,ProductNode_POSIT15Output_18);

ProductNode_POSIT16: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT16weight,ProductNode_POSIT15Output_18,ProductNode_POSIT16Output_19);

ProductNode_POSIT17: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT17weight,vb8,ProductNode_POSIT17Output_20);

ProductNode_POSIT18: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT18weight,ProductNode_POSIT17Output_20,ProductNode_POSIT18Output_21);

SumNode_POSIT3: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT18Output_21,ProductNode_POSIT16Output_19,SumNode_POSIT3Output_22);

ProductNode_POSIT19: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT3Output_22,ProductNode_POSIT14Output_17,ProductNode_POSIT19Output_23);

SumNode_POSIT4: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT19Output_23,ProductNode_POSIT11Output_13,SumNode_POSIT4Output_24);

ProductNode_POSIT20: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT4Output_24,ProductNode_POSIT3Output_3,ProductNode_POSIT20Output_25);

ProductNode_POSIT21: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT21weight,vb2,ProductNode_POSIT21Output_26);

ProductNode_POSIT25: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT25weight,v8,ProductNode_POSIT25Output_31);

ProductNode_POSIT26: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT26weight,ProductNode_POSIT25Output_31,ProductNode_POSIT26Output_32);

ProductNode_POSIT27: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT27weight,vb8,ProductNode_POSIT27Output_33);

ProductNode_POSIT28: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT28weight,ProductNode_POSIT27Output_33,ProductNode_POSIT28Output_34);

SumNode_POSIT6: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT28Output_34,ProductNode_POSIT26Output_32,SumNode_POSIT6Output_35);

ProductNode_POSIT29: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT6Output_35,ProductNode_POSIT6Output_7,ProductNode_POSIT29Output_36);

ProductNode_POSIT33: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT33weight,v8,ProductNode_POSIT33Output_41);

ProductNode_POSIT34: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT34weight,ProductNode_POSIT33Output_41,ProductNode_POSIT34Output_42);

ProductNode_POSIT35: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT35weight,vb8,ProductNode_POSIT35Output_43);

ProductNode_POSIT36: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT36weight,ProductNode_POSIT35Output_43,ProductNode_POSIT36Output_44);

SumNode_POSIT8: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT36Output_44,ProductNode_POSIT34Output_42,SumNode_POSIT8Output_45);

ProductNode_POSIT37: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT8Output_45,ProductNode_POSIT14Output_17,ProductNode_POSIT37Output_46);

SumNode_POSIT9: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT37Output_46,ProductNode_POSIT29Output_36,SumNode_POSIT9Output_47);

ProductNode_POSIT38: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT9Output_47,ProductNode_POSIT21Output_26,ProductNode_POSIT38Output_48);

SumNode_POSIT10: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT38Output_48,ProductNode_POSIT20Output_25,SumNode_POSIT10Output_49);

ProductNode_POSIT39: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT10Output_49,ProductNode_POSIT2Output_2,ProductNode_POSIT39Output_50);

ProductNode_POSIT40: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT40weight,v10,ProductNode_POSIT40Output_51);

ProductNode_POSIT41: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT41weight,v5,ProductNode_POSIT41Output_52);

ProductNode_POSIT42: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT42weight,ProductNode_POSIT41Output_52,ProductNode_POSIT42Output_53);

ProductNode_POSIT43: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT43weight,ProductNode_POSIT42Output_53,ProductNode_POSIT43Output_54);

ProductNode_POSIT44: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT44weight,ProductNode_POSIT43Output_54,ProductNode_POSIT44Output_55);

ProductNode_POSIT45: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT45weight,vb5,ProductNode_POSIT45Output_56);

ProductNode_POSIT46: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT46weight,ProductNode_POSIT45Output_56,ProductNode_POSIT46Output_57);

ProductNode_POSIT47: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT47weight,ProductNode_POSIT46Output_57,ProductNode_POSIT47Output_58);

ProductNode_POSIT48: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT48weight,ProductNode_POSIT47Output_58,ProductNode_POSIT48Output_59);

SumNode_POSIT11: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT48Output_59,ProductNode_POSIT44Output_55,SumNode_POSIT11Output_60);

ProductNode_POSIT49: entity work.PositMult_23_6_comb_uid2(arch)
port map(v16,SumNode_POSIT11Output_60,ProductNode_POSIT49Output_61);

ProductNode_POSIT50: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT50weight,ProductNode_POSIT49Output_61,ProductNode_POSIT50Output_62);

ProductNode_POSIT53: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT53weight,ProductNode_POSIT42Output_53,ProductNode_POSIT53Output_65);

ProductNode_POSIT54: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT54weight,ProductNode_POSIT53Output_65,ProductNode_POSIT54Output_66);

ProductNode_POSIT57: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT57weight,ProductNode_POSIT46Output_57,ProductNode_POSIT57Output_69);

ProductNode_POSIT58: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT58weight,ProductNode_POSIT57Output_69,ProductNode_POSIT58Output_70);

SumNode_POSIT12: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT58Output_70,ProductNode_POSIT54Output_66,SumNode_POSIT12Output_71);

ProductNode_POSIT59: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb16,SumNode_POSIT12Output_71,ProductNode_POSIT59Output_72);

ProductNode_POSIT60: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT60weight,ProductNode_POSIT59Output_72,ProductNode_POSIT60Output_73);

SumNode_POSIT13: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT60Output_73,ProductNode_POSIT50Output_62,SumNode_POSIT13Output_74);

ProductNode_POSIT61: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT13Output_74,ProductNode_POSIT40Output_51,ProductNode_POSIT61Output_75);

ProductNode_POSIT62: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT62weight,ProductNode_POSIT61Output_75,ProductNode_POSIT62Output_76);

ProductNode_POSIT63: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT63weight,v14,ProductNode_POSIT63Output_77);

ProductNode_POSIT64: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT64weight,vb14,ProductNode_POSIT64Output_78);

SumNode_POSIT14: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT64Output_78,ProductNode_POSIT63Output_77,SumNode_POSIT14Output_79);

ProductNode_POSIT65: entity work.PositMult_23_6_comb_uid2(arch)
port map(v15,SumNode_POSIT14Output_79,ProductNode_POSIT65Output_80);

ProductNode_POSIT66: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT66weight,ProductNode_POSIT65Output_80,ProductNode_POSIT66Output_81);

ProductNode_POSIT67: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT67weight,v14,ProductNode_POSIT67Output_82);

ProductNode_POSIT68: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT68weight,vb14,ProductNode_POSIT68Output_83);

SumNode_POSIT15: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT68Output_83,ProductNode_POSIT67Output_82,SumNode_POSIT15Output_84);

ProductNode_POSIT69: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb15,SumNode_POSIT15Output_84,ProductNode_POSIT69Output_85);

ProductNode_POSIT70: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT70weight,ProductNode_POSIT69Output_85,ProductNode_POSIT70Output_86);

SumNode_POSIT16: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT70Output_86,ProductNode_POSIT66Output_81,SumNode_POSIT16Output_87);

ProductNode_POSIT71: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT16Output_87,ProductNode_POSIT62Output_76,ProductNode_POSIT71Output_88);

ProductNode_POSIT72: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT72weight,vb10,ProductNode_POSIT72Output_89);

ProductNode_POSIT73: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT73weight,v5,ProductNode_POSIT73Output_90);

ProductNode_POSIT74: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT74weight,ProductNode_POSIT73Output_90,ProductNode_POSIT74Output_91);

ProductNode_POSIT75: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT75weight,ProductNode_POSIT74Output_91,ProductNode_POSIT75Output_92);

ProductNode_POSIT76: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT76weight,ProductNode_POSIT75Output_92,ProductNode_POSIT76Output_93);

ProductNode_POSIT77: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT77weight,vb5,ProductNode_POSIT77Output_94);

ProductNode_POSIT78: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT78weight,ProductNode_POSIT77Output_94,ProductNode_POSIT78Output_95);

ProductNode_POSIT79: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT79weight,ProductNode_POSIT78Output_95,ProductNode_POSIT79Output_96);

ProductNode_POSIT80: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT80weight,ProductNode_POSIT79Output_96,ProductNode_POSIT80Output_97);

SumNode_POSIT17: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT80Output_97,ProductNode_POSIT76Output_93,SumNode_POSIT17Output_98);

ProductNode_POSIT81: entity work.PositMult_23_6_comb_uid2(arch)
port map(v16,SumNode_POSIT17Output_98,ProductNode_POSIT81Output_99);

ProductNode_POSIT82: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT82weight,ProductNode_POSIT81Output_99,ProductNode_POSIT82Output_100);

ProductNode_POSIT85: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT85weight,ProductNode_POSIT74Output_91,ProductNode_POSIT85Output_103);

ProductNode_POSIT86: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT86weight,ProductNode_POSIT85Output_103,ProductNode_POSIT86Output_104);

ProductNode_POSIT89: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT89weight,ProductNode_POSIT78Output_95,ProductNode_POSIT89Output_107);

ProductNode_POSIT90: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT90weight,ProductNode_POSIT89Output_107,ProductNode_POSIT90Output_108);

SumNode_POSIT18: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT90Output_108,ProductNode_POSIT86Output_104,SumNode_POSIT18Output_109);

ProductNode_POSIT91: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb16,SumNode_POSIT18Output_109,ProductNode_POSIT91Output_110);

ProductNode_POSIT92: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT92weight,ProductNode_POSIT91Output_110,ProductNode_POSIT92Output_111);

SumNode_POSIT19: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT92Output_111,ProductNode_POSIT82Output_100,SumNode_POSIT19Output_112);

ProductNode_POSIT93: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT19Output_112,ProductNode_POSIT72Output_89,ProductNode_POSIT93Output_113);

ProductNode_POSIT94: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT94weight,ProductNode_POSIT93Output_113,ProductNode_POSIT94Output_114);

ProductNode_POSIT98: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT98weight,ProductNode_POSIT65Output_80,ProductNode_POSIT98Output_119);

ProductNode_POSIT102: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT102weight,ProductNode_POSIT69Output_85,ProductNode_POSIT102Output_124);

SumNode_POSIT22: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT102Output_124,ProductNode_POSIT98Output_119,SumNode_POSIT22Output_125);

ProductNode_POSIT103: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT22Output_125,ProductNode_POSIT94Output_114,ProductNode_POSIT103Output_126);

SumNode_POSIT23: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT103Output_126,ProductNode_POSIT71Output_88,SumNode_POSIT23Output_127);

ProductNode_POSIT104: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT23Output_127,ProductNode_POSIT39Output_50,ProductNode_POSIT104Output_128);

ProductNode_POSIT105: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT105weight,vb11,ProductNode_POSIT105Output_129);

ProductNode_POSIT106: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT106weight,ProductNode_POSIT105Output_129,ProductNode_POSIT106Output_130);

ProductNode_POSIT112: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT112weight,ProductNode_POSIT7Output_8,ProductNode_POSIT112Output_137);

ProductNode_POSIT114: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT114weight,ProductNode_POSIT9Output_10,ProductNode_POSIT114Output_139);

SumNode_POSIT25: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT114Output_139,ProductNode_POSIT112Output_137,SumNode_POSIT25Output_140);

ProductNode_POSIT115: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT25Output_140,ProductNode_POSIT6Output_7,ProductNode_POSIT115Output_141);

ProductNode_POSIT120: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT120weight,ProductNode_POSIT15Output_18,ProductNode_POSIT120Output_147);

ProductNode_POSIT122: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT122weight,ProductNode_POSIT17Output_20,ProductNode_POSIT122Output_149);

SumNode_POSIT27: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT122Output_149,ProductNode_POSIT120Output_147,SumNode_POSIT27Output_150);

ProductNode_POSIT123: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT27Output_150,ProductNode_POSIT14Output_17,ProductNode_POSIT123Output_151);

SumNode_POSIT28: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT123Output_151,ProductNode_POSIT115Output_141,SumNode_POSIT28Output_152);

ProductNode_POSIT124: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT28Output_152,ProductNode_POSIT3Output_3,ProductNode_POSIT124Output_153);

ProductNode_POSIT130: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT130weight,ProductNode_POSIT25Output_31,ProductNode_POSIT130Output_160);

ProductNode_POSIT132: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT132weight,ProductNode_POSIT27Output_33,ProductNode_POSIT132Output_162);

SumNode_POSIT30: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT132Output_162,ProductNode_POSIT130Output_160,SumNode_POSIT30Output_163);

ProductNode_POSIT133: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT30Output_163,ProductNode_POSIT6Output_7,ProductNode_POSIT133Output_164);

ProductNode_POSIT138: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT138weight,ProductNode_POSIT33Output_41,ProductNode_POSIT138Output_170);

ProductNode_POSIT140: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT140weight,ProductNode_POSIT35Output_43,ProductNode_POSIT140Output_172);

SumNode_POSIT32: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT140Output_172,ProductNode_POSIT138Output_170,SumNode_POSIT32Output_173);

ProductNode_POSIT141: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT32Output_173,ProductNode_POSIT14Output_17,ProductNode_POSIT141Output_174);

SumNode_POSIT33: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT141Output_174,ProductNode_POSIT133Output_164,SumNode_POSIT33Output_175);

ProductNode_POSIT142: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT33Output_175,ProductNode_POSIT21Output_26,ProductNode_POSIT142Output_176);

SumNode_POSIT34: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT142Output_176,ProductNode_POSIT124Output_153,SumNode_POSIT34Output_177);

ProductNode_POSIT143: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT34Output_177,ProductNode_POSIT106Output_130,ProductNode_POSIT143Output_178);

ProductNode_POSIT166: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT166weight,ProductNode_POSIT61Output_75,ProductNode_POSIT166Output_204);

ProductNode_POSIT170: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT170weight,ProductNode_POSIT65Output_80,ProductNode_POSIT170Output_209);

ProductNode_POSIT174: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT174weight,ProductNode_POSIT69Output_85,ProductNode_POSIT174Output_214);

SumNode_POSIT40: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT174Output_214,ProductNode_POSIT170Output_209,SumNode_POSIT40Output_215);

ProductNode_POSIT175: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT40Output_215,ProductNode_POSIT166Output_204,ProductNode_POSIT175Output_216);

ProductNode_POSIT198: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT198weight,ProductNode_POSIT93Output_113,ProductNode_POSIT198Output_242);

ProductNode_POSIT202: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT202weight,ProductNode_POSIT65Output_80,ProductNode_POSIT202Output_247);

ProductNode_POSIT206: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT206weight,ProductNode_POSIT69Output_85,ProductNode_POSIT206Output_252);

SumNode_POSIT46: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT206Output_252,ProductNode_POSIT202Output_247,SumNode_POSIT46Output_253);

ProductNode_POSIT207: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT46Output_253,ProductNode_POSIT198Output_242,ProductNode_POSIT207Output_254);

SumNode_POSIT47: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT207Output_254,ProductNode_POSIT175Output_216,SumNode_POSIT47Output_255);

ProductNode_POSIT208: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT47Output_255,ProductNode_POSIT143Output_178,ProductNode_POSIT208Output_256);

SumNode_POSIT48: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT208Output_256,ProductNode_POSIT104Output_128,SumNode_POSIT48Output_257);

ProductNode_POSIT209: entity work.PositMult_23_6_comb_uid2(arch)
port map(v13,SumNode_POSIT48Output_257,ProductNode_POSIT209Output_258);

ProductNode_POSIT211: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT211weight,ProductNode_POSIT1Output_1,ProductNode_POSIT211Output_260);

ProductNode_POSIT248: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT59Output_307,ProductNode_POSIT211Output_260,ProductNode_POSIT248Output_308);

ProductNode_POSIT272: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT272weight,v14,ProductNode_POSIT272Output_335);

ProductNode_POSIT273: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT273weight,vb14,ProductNode_POSIT273Output_336);

SumNode_POSIT63: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT273Output_336,ProductNode_POSIT272Output_335,SumNode_POSIT63Output_337);

ProductNode_POSIT274: entity work.PositMult_23_6_comb_uid2(arch)
port map(v15,SumNode_POSIT63Output_337,ProductNode_POSIT274Output_338);

ProductNode_POSIT275: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT275weight,ProductNode_POSIT274Output_338,ProductNode_POSIT275Output_339);

ProductNode_POSIT276: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT276weight,v14,ProductNode_POSIT276Output_340);

ProductNode_POSIT277: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT277weight,vb14,ProductNode_POSIT277Output_341);

SumNode_POSIT64: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT277Output_341,ProductNode_POSIT276Output_340,SumNode_POSIT64Output_342);

ProductNode_POSIT278: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb15,SumNode_POSIT64Output_342,ProductNode_POSIT278Output_343);

ProductNode_POSIT279: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT279weight,ProductNode_POSIT278Output_343,ProductNode_POSIT279Output_344);

SumNode_POSIT65: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT279Output_344,ProductNode_POSIT275Output_339,SumNode_POSIT65Output_345);

ProductNode_POSIT280: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT65Output_345,ProductNode_POSIT62Output_76,ProductNode_POSIT280Output_346);

ProductNode_POSIT307: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT307weight,ProductNode_POSIT274Output_338,ProductNode_POSIT307Output_377);

ProductNode_POSIT311: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT311weight,ProductNode_POSIT278Output_343,ProductNode_POSIT311Output_382);

SumNode_POSIT71: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT311Output_382,ProductNode_POSIT307Output_377,SumNode_POSIT71Output_383);

ProductNode_POSIT312: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT71Output_383,ProductNode_POSIT94Output_114,ProductNode_POSIT312Output_384);

SumNode_POSIT72: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT312Output_384,ProductNode_POSIT280Output_346,SumNode_POSIT72Output_385);

ProductNode_POSIT313: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT72Output_385,ProductNode_POSIT248Output_308,ProductNode_POSIT313Output_386);

ProductNode_POSIT315: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT315weight,ProductNode_POSIT105Output_129,ProductNode_POSIT315Output_388);

ProductNode_POSIT352: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT83Output_435,ProductNode_POSIT315Output_388,ProductNode_POSIT352Output_436);

ProductNode_POSIT379: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT379weight,ProductNode_POSIT274Output_338,ProductNode_POSIT379Output_467);

ProductNode_POSIT383: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT383weight,ProductNode_POSIT278Output_343,ProductNode_POSIT383Output_472);

SumNode_POSIT89: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT383Output_472,ProductNode_POSIT379Output_467,SumNode_POSIT89Output_473);

ProductNode_POSIT384: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT89Output_473,ProductNode_POSIT166Output_204,ProductNode_POSIT384Output_474);

ProductNode_POSIT411: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT411weight,ProductNode_POSIT274Output_338,ProductNode_POSIT411Output_505);

ProductNode_POSIT415: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT415weight,ProductNode_POSIT278Output_343,ProductNode_POSIT415Output_510);

SumNode_POSIT95: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT415Output_510,ProductNode_POSIT411Output_505,SumNode_POSIT95Output_511);

ProductNode_POSIT416: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT95Output_511,ProductNode_POSIT198Output_242,ProductNode_POSIT416Output_512);

SumNode_POSIT96: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT416Output_512,ProductNode_POSIT384Output_474,SumNode_POSIT96Output_513);

ProductNode_POSIT417: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT96Output_513,ProductNode_POSIT352Output_436,ProductNode_POSIT417Output_514);

SumNode_POSIT97: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT417Output_514,ProductNode_POSIT313Output_386,SumNode_POSIT97Output_515);

ProductNode_POSIT418: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb13,SumNode_POSIT97Output_515,ProductNode_POSIT418Output_516);

SumNode_POSIT98: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT418Output_516,ProductNode_POSIT209Output_258,SumNode_POSIT98Output_517);

ProductNode_POSIT419: entity work.PositMult_23_6_comb_uid2(arch)
port map(v3,SumNode_POSIT98Output_517,ProductNode_POSIT419Output_518);

ProductNode_POSIT422: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT422weight,v2,ProductNode_POSIT422Output_521);

ProductNode_POSIT439: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT103Output_542,ProductNode_POSIT422Output_521,ProductNode_POSIT439Output_543);

ProductNode_POSIT440: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT440weight,vb2,ProductNode_POSIT440Output_544);

ProductNode_POSIT457: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT108Output_565,ProductNode_POSIT440Output_544,ProductNode_POSIT457Output_566);

SumNode_POSIT109: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT457Output_566,ProductNode_POSIT439Output_543,SumNode_POSIT109Output_567);

ProductNode_POSIT458: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT109Output_567,ProductNode_POSIT2Output_2,ProductNode_POSIT458Output_568);

ProductNode_POSIT463: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT463weight,ProductNode_POSIT43Output_54,ProductNode_POSIT463Output_573);

ProductNode_POSIT467: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT467weight,ProductNode_POSIT47Output_58,ProductNode_POSIT467Output_577);

SumNode_POSIT110: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT467Output_577,ProductNode_POSIT463Output_573,SumNode_POSIT110Output_578);

ProductNode_POSIT468: entity work.PositMult_23_6_comb_uid2(arch)
port map(v16,SumNode_POSIT110Output_578,ProductNode_POSIT468Output_579);

ProductNode_POSIT469: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT469weight,ProductNode_POSIT468Output_579,ProductNode_POSIT469Output_580);

ProductNode_POSIT473: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT473weight,ProductNode_POSIT53Output_65,ProductNode_POSIT473Output_584);

ProductNode_POSIT477: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT477weight,ProductNode_POSIT57Output_69,ProductNode_POSIT477Output_588);

SumNode_POSIT111: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT477Output_588,ProductNode_POSIT473Output_584,SumNode_POSIT111Output_589);

ProductNode_POSIT478: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb16,SumNode_POSIT111Output_589,ProductNode_POSIT478Output_590);

ProductNode_POSIT479: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT479weight,ProductNode_POSIT478Output_590,ProductNode_POSIT479Output_591);

SumNode_POSIT112: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT479Output_591,ProductNode_POSIT469Output_580,SumNode_POSIT112Output_592);

ProductNode_POSIT480: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT112Output_592,ProductNode_POSIT40Output_51,ProductNode_POSIT480Output_593);

ProductNode_POSIT481: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT481weight,ProductNode_POSIT480Output_593,ProductNode_POSIT481Output_594);

ProductNode_POSIT485: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT485weight,ProductNode_POSIT65Output_80,ProductNode_POSIT485Output_599);

ProductNode_POSIT489: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT489weight,ProductNode_POSIT69Output_85,ProductNode_POSIT489Output_604);

SumNode_POSIT115: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT489Output_604,ProductNode_POSIT485Output_599,SumNode_POSIT115Output_605);

ProductNode_POSIT490: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT115Output_605,ProductNode_POSIT481Output_594,ProductNode_POSIT490Output_606);

ProductNode_POSIT495: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT495weight,ProductNode_POSIT75Output_92,ProductNode_POSIT495Output_611);

ProductNode_POSIT499: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT499weight,ProductNode_POSIT79Output_96,ProductNode_POSIT499Output_615);

SumNode_POSIT116: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT499Output_615,ProductNode_POSIT495Output_611,SumNode_POSIT116Output_616);

ProductNode_POSIT500: entity work.PositMult_23_6_comb_uid2(arch)
port map(v16,SumNode_POSIT116Output_616,ProductNode_POSIT500Output_617);

ProductNode_POSIT501: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT501weight,ProductNode_POSIT500Output_617,ProductNode_POSIT501Output_618);

ProductNode_POSIT505: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT505weight,ProductNode_POSIT85Output_103,ProductNode_POSIT505Output_622);

SumNode_POSIT117: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT509Output_626,ProductNode_POSIT505Output_622,SumNode_POSIT117Output_627);

ProductNode_POSIT510: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb16,SumNode_POSIT117Output_627,ProductNode_POSIT510Output_628);

ProductNode_POSIT511: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT511weight,ProductNode_POSIT510Output_628,ProductNode_POSIT511Output_629);

SumNode_POSIT118: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT511Output_629,ProductNode_POSIT501Output_618,SumNode_POSIT118Output_630);

ProductNode_POSIT512: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT118Output_630,ProductNode_POSIT72Output_89,ProductNode_POSIT512Output_631);

ProductNode_POSIT513: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT513weight,ProductNode_POSIT512Output_631,ProductNode_POSIT513Output_632);

ProductNode_POSIT517: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT517weight,ProductNode_POSIT65Output_80,ProductNode_POSIT517Output_637);

ProductNode_POSIT521: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT521weight,ProductNode_POSIT69Output_85,ProductNode_POSIT521Output_642);

SumNode_POSIT121: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT521Output_642,ProductNode_POSIT517Output_637,SumNode_POSIT121Output_643);

ProductNode_POSIT522: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT121Output_643,ProductNode_POSIT513Output_632,ProductNode_POSIT522Output_644);

SumNode_POSIT122: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT522Output_644,ProductNode_POSIT490Output_606,SumNode_POSIT122Output_645);

ProductNode_POSIT523: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT122Output_645,ProductNode_POSIT458Output_568,ProductNode_POSIT523Output_646);

ProductNode_POSIT543: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT28Output_152,ProductNode_POSIT422Output_521,ProductNode_POSIT543Output_671);

ProductNode_POSIT561: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT33Output_175,ProductNode_POSIT440Output_544,ProductNode_POSIT561Output_694);

SumNode_POSIT133: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT561Output_694,ProductNode_POSIT543Output_671,SumNode_POSIT133Output_695);

ProductNode_POSIT562: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT133Output_695,ProductNode_POSIT106Output_130,ProductNode_POSIT562Output_696);

ProductNode_POSIT585: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT585weight,ProductNode_POSIT480Output_593,ProductNode_POSIT585Output_722);

ProductNode_POSIT589: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT589weight,ProductNode_POSIT65Output_80,ProductNode_POSIT589Output_727);

ProductNode_POSIT593: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT593weight,ProductNode_POSIT69Output_85,ProductNode_POSIT593Output_732);

SumNode_POSIT139: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT593Output_732,ProductNode_POSIT589Output_727,SumNode_POSIT139Output_733);

ProductNode_POSIT594: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT139Output_733,ProductNode_POSIT585Output_722,ProductNode_POSIT594Output_734);

ProductNode_POSIT617: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT617weight,ProductNode_POSIT512Output_631,ProductNode_POSIT617Output_760);

ProductNode_POSIT621: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT621weight,ProductNode_POSIT65Output_80,ProductNode_POSIT621Output_765);

ProductNode_POSIT625: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT625weight,ProductNode_POSIT69Output_85,ProductNode_POSIT625Output_770);

SumNode_POSIT145: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT625Output_770,ProductNode_POSIT621Output_765,SumNode_POSIT145Output_771);

ProductNode_POSIT626: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT145Output_771,ProductNode_POSIT617Output_760,ProductNode_POSIT626Output_772);

SumNode_POSIT146: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT626Output_772,ProductNode_POSIT594Output_734,SumNode_POSIT146Output_773);

ProductNode_POSIT627: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT146Output_773,ProductNode_POSIT562Output_696,ProductNode_POSIT627Output_774);

SumNode_POSIT147: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT627Output_774,ProductNode_POSIT523Output_646,SumNode_POSIT147Output_775);

ProductNode_POSIT628: entity work.PositMult_23_6_comb_uid2(arch)
port map(v13,SumNode_POSIT147Output_775,ProductNode_POSIT628Output_776);

ProductNode_POSIT667: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT158Output_825,ProductNode_POSIT211Output_260,ProductNode_POSIT667Output_826);

ProductNode_POSIT694: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT694weight,ProductNode_POSIT274Output_338,ProductNode_POSIT694Output_857);

ProductNode_POSIT698: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT698weight,ProductNode_POSIT278Output_343,ProductNode_POSIT698Output_862);

SumNode_POSIT164: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT698Output_862,ProductNode_POSIT694Output_857,SumNode_POSIT164Output_863);

ProductNode_POSIT699: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT164Output_863,ProductNode_POSIT481Output_594,ProductNode_POSIT699Output_864);

ProductNode_POSIT726: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT726weight,ProductNode_POSIT274Output_338,ProductNode_POSIT726Output_895);

ProductNode_POSIT730: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT730weight,ProductNode_POSIT278Output_343,ProductNode_POSIT730Output_900);

SumNode_POSIT170: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT730Output_900,ProductNode_POSIT726Output_895,SumNode_POSIT170Output_901);

ProductNode_POSIT731: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT170Output_901,ProductNode_POSIT513Output_632,ProductNode_POSIT731Output_902);

SumNode_POSIT171: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT731Output_902,ProductNode_POSIT699Output_864,SumNode_POSIT171Output_903);

ProductNode_POSIT732: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT171Output_903,ProductNode_POSIT667Output_826,ProductNode_POSIT732Output_904);

ProductNode_POSIT771: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT182Output_953,ProductNode_POSIT315Output_388,ProductNode_POSIT771Output_954);

ProductNode_POSIT798: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT798weight,ProductNode_POSIT274Output_338,ProductNode_POSIT798Output_985);

ProductNode_POSIT802: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT802weight,ProductNode_POSIT278Output_343,ProductNode_POSIT802Output_990);

SumNode_POSIT188: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT802Output_990,ProductNode_POSIT798Output_985,SumNode_POSIT188Output_991);

ProductNode_POSIT803: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT188Output_991,ProductNode_POSIT585Output_722,ProductNode_POSIT803Output_992);

ProductNode_POSIT830: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT830weight,ProductNode_POSIT274Output_338,ProductNode_POSIT830Output_1023);

ProductNode_POSIT834: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT834weight,ProductNode_POSIT278Output_343,ProductNode_POSIT834Output_1028);

SumNode_POSIT194: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT834Output_1028,ProductNode_POSIT830Output_1023,SumNode_POSIT194Output_1029);

ProductNode_POSIT835: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT194Output_1029,ProductNode_POSIT617Output_760,ProductNode_POSIT835Output_1030);

SumNode_POSIT195: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT835Output_1030,ProductNode_POSIT803Output_992,SumNode_POSIT195Output_1031);

ProductNode_POSIT836: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT195Output_1031,ProductNode_POSIT771Output_954,ProductNode_POSIT836Output_1032);

SumNode_POSIT196: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT836Output_1032,ProductNode_POSIT732Output_904,SumNode_POSIT196Output_1033);

ProductNode_POSIT837: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb13,SumNode_POSIT196Output_1033,ProductNode_POSIT837Output_1034);

SumNode_POSIT197: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT837Output_1034,ProductNode_POSIT628Output_776,SumNode_POSIT197Output_1035);

ProductNode_POSIT838: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb3,SumNode_POSIT197Output_1035,ProductNode_POSIT838Output_1036);

SumNode_POSIT198: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT838Output_1036,ProductNode_POSIT419Output_518,SumNode_POSIT198Output_1037);

ProductNode_POSIT839: entity work.PositMult_23_6_comb_uid2(arch)
port map(v4,SumNode_POSIT198Output_1037,ProductNode_POSIT839Output_1038);

ProductNode_POSIT840: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT840weight,v11,ProductNode_POSIT840Output_1039);

ProductNode_POSIT841: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT841weight,ProductNode_POSIT840Output_1039,ProductNode_POSIT841Output_1040);

ProductNode_POSIT842: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT842weight,v2,ProductNode_POSIT842Output_1041);

ProductNode_POSIT843: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT843weight,v7,ProductNode_POSIT843Output_1042);

ProductNode_POSIT844: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT844weight,vb7,ProductNode_POSIT844Output_1043);

SumNode_POSIT199: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT844Output_1043,ProductNode_POSIT843Output_1042,SumNode_POSIT199Output_1044);

ProductNode_POSIT845: entity work.PositMult_23_6_comb_uid2(arch)
port map(v1,SumNode_POSIT199Output_1044,ProductNode_POSIT845Output_1045);

ProductNode_POSIT850: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT200Output_1050,ProductNode_POSIT845Output_1045,ProductNode_POSIT850Output_1051);

ProductNode_POSIT851: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT851weight,v7,ProductNode_POSIT851Output_1052);

ProductNode_POSIT852: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT852weight,vb7,ProductNode_POSIT852Output_1053);

SumNode_POSIT201: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT852Output_1053,ProductNode_POSIT851Output_1052,SumNode_POSIT201Output_1054);

ProductNode_POSIT853: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb1,SumNode_POSIT201Output_1054,ProductNode_POSIT853Output_1055);

ProductNode_POSIT858: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT202Output_1060,ProductNode_POSIT853Output_1055,ProductNode_POSIT858Output_1061);

SumNode_POSIT203: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT858Output_1061,ProductNode_POSIT850Output_1051,SumNode_POSIT203Output_1062);

ProductNode_POSIT859: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT203Output_1062,ProductNode_POSIT842Output_1041,ProductNode_POSIT859Output_1063);

ProductNode_POSIT860: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT860weight,vb2,ProductNode_POSIT860Output_1064);

ProductNode_POSIT868: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT6Output_35,ProductNode_POSIT845Output_1045,ProductNode_POSIT868Output_1074);

ProductNode_POSIT876: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT8Output_45,ProductNode_POSIT853Output_1055,ProductNode_POSIT876Output_1084);

SumNode_POSIT208: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT876Output_1084,ProductNode_POSIT868Output_1074,SumNode_POSIT208Output_1085);

ProductNode_POSIT877: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT208Output_1085,ProductNode_POSIT860Output_1064,ProductNode_POSIT877Output_1086);

SumNode_POSIT209: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT877Output_1086,ProductNode_POSIT859Output_1063,SumNode_POSIT209Output_1087);

ProductNode_POSIT878: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT209Output_1087,ProductNode_POSIT841Output_1040,ProductNode_POSIT878Output_1088);

ProductNode_POSIT889: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT889weight,ProductNode_POSIT49Output_61,ProductNode_POSIT889Output_1100);

ProductNode_POSIT899: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT899weight,ProductNode_POSIT59Output_72,ProductNode_POSIT899Output_1111);

SumNode_POSIT212: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT899Output_1111,ProductNode_POSIT889Output_1100,SumNode_POSIT212Output_1112);

ProductNode_POSIT900: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT212Output_1112,ProductNode_POSIT40Output_51,ProductNode_POSIT900Output_1113);

ProductNode_POSIT901: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT901weight,ProductNode_POSIT900Output_1113,ProductNode_POSIT901Output_1114);

ProductNode_POSIT902: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT902weight,v14,ProductNode_POSIT902Output_1115);

ProductNode_POSIT903: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT903weight,vb14,ProductNode_POSIT903Output_1116);

SumNode_POSIT213: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT903Output_1116,ProductNode_POSIT902Output_1115,SumNode_POSIT213Output_1117);

ProductNode_POSIT904: entity work.PositMult_23_6_comb_uid2(arch)
port map(v15,SumNode_POSIT213Output_1117,ProductNode_POSIT904Output_1118);

ProductNode_POSIT905: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT905weight,ProductNode_POSIT904Output_1118,ProductNode_POSIT905Output_1119);

ProductNode_POSIT906: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT906weight,v14,ProductNode_POSIT906Output_1120);

ProductNode_POSIT907: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT907weight,vb14,ProductNode_POSIT907Output_1121);

SumNode_POSIT214: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT907Output_1121,ProductNode_POSIT906Output_1120,SumNode_POSIT214Output_1122);

ProductNode_POSIT908: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb15,SumNode_POSIT214Output_1122,ProductNode_POSIT908Output_1123);

ProductNode_POSIT909: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT909weight,ProductNode_POSIT908Output_1123,ProductNode_POSIT909Output_1124);

SumNode_POSIT215: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT909Output_1124,ProductNode_POSIT905Output_1119,SumNode_POSIT215Output_1125);

ProductNode_POSIT910: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT215Output_1125,ProductNode_POSIT901Output_1114,ProductNode_POSIT910Output_1126);

ProductNode_POSIT921: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT921weight,ProductNode_POSIT81Output_99,ProductNode_POSIT921Output_1138);

ProductNode_POSIT931: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT931weight,ProductNode_POSIT91Output_110,ProductNode_POSIT931Output_1149);

SumNode_POSIT218: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT931Output_1149,ProductNode_POSIT921Output_1138,SumNode_POSIT218Output_1150);

ProductNode_POSIT932: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT218Output_1150,ProductNode_POSIT72Output_89,ProductNode_POSIT932Output_1151);

ProductNode_POSIT933: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT933weight,ProductNode_POSIT932Output_1151,ProductNode_POSIT933Output_1152);

ProductNode_POSIT937: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT937weight,ProductNode_POSIT904Output_1118,ProductNode_POSIT937Output_1157);

ProductNode_POSIT941: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT941weight,ProductNode_POSIT908Output_1123,ProductNode_POSIT941Output_1162);

SumNode_POSIT221: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT941Output_1162,ProductNode_POSIT937Output_1157,SumNode_POSIT221Output_1163);

ProductNode_POSIT942: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT221Output_1163,ProductNode_POSIT933Output_1152,ProductNode_POSIT942Output_1164);

SumNode_POSIT222: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT942Output_1164,ProductNode_POSIT910Output_1126,SumNode_POSIT222Output_1165);

ProductNode_POSIT943: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT222Output_1165,ProductNode_POSIT878Output_1088,ProductNode_POSIT943Output_1166);

ProductNode_POSIT944: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT944weight,vb11,ProductNode_POSIT944Output_1167);

ProductNode_POSIT945: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT945weight,ProductNode_POSIT944Output_1167,ProductNode_POSIT945Output_1168);

ProductNode_POSIT954: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT25Output_140,ProductNode_POSIT845Output_1045,ProductNode_POSIT954Output_1179);

ProductNode_POSIT962: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT27Output_150,ProductNode_POSIT853Output_1055,ProductNode_POSIT962Output_1189);

SumNode_POSIT227: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT962Output_1189,ProductNode_POSIT954Output_1179,SumNode_POSIT227Output_1190);

ProductNode_POSIT963: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT227Output_1190,ProductNode_POSIT842Output_1041,ProductNode_POSIT963Output_1191);

ProductNode_POSIT972: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT30Output_163,ProductNode_POSIT845Output_1045,ProductNode_POSIT972Output_1202);

ProductNode_POSIT980: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT32Output_173,ProductNode_POSIT853Output_1055,ProductNode_POSIT980Output_1212);

SumNode_POSIT232: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT980Output_1212,ProductNode_POSIT972Output_1202,SumNode_POSIT232Output_1213);

ProductNode_POSIT981: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT232Output_1213,ProductNode_POSIT860Output_1064,ProductNode_POSIT981Output_1214);

SumNode_POSIT233: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT981Output_1214,ProductNode_POSIT963Output_1191,SumNode_POSIT233Output_1215);

ProductNode_POSIT982: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT233Output_1215,ProductNode_POSIT945Output_1168,ProductNode_POSIT982Output_1216);

ProductNode_POSIT1005: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1005weight,ProductNode_POSIT900Output_1113,ProductNode_POSIT1005Output_1242);

ProductNode_POSIT1009: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1009weight,ProductNode_POSIT904Output_1118,ProductNode_POSIT1009Output_1247);

ProductNode_POSIT1013: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1013weight,ProductNode_POSIT908Output_1123,ProductNode_POSIT1013Output_1252);

SumNode_POSIT239: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT1013Output_1252,ProductNode_POSIT1009Output_1247,SumNode_POSIT239Output_1253);

ProductNode_POSIT1014: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT239Output_1253,ProductNode_POSIT1005Output_1242,ProductNode_POSIT1014Output_1254);

ProductNode_POSIT1037: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1037weight,ProductNode_POSIT932Output_1151,ProductNode_POSIT1037Output_1280);

ProductNode_POSIT1041: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1041weight,ProductNode_POSIT904Output_1118,ProductNode_POSIT1041Output_1285);

ProductNode_POSIT1045: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1045weight,ProductNode_POSIT908Output_1123,ProductNode_POSIT1045Output_1290);

SumNode_POSIT245: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT1045Output_1290,ProductNode_POSIT1041Output_1285,SumNode_POSIT245Output_1291);

ProductNode_POSIT1046: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT245Output_1291,ProductNode_POSIT1037Output_1280,ProductNode_POSIT1046Output_1292);

SumNode_POSIT246: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT1046Output_1292,ProductNode_POSIT1014Output_1254,SumNode_POSIT246Output_1293);

ProductNode_POSIT1047: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT246Output_1293,ProductNode_POSIT982Output_1216,ProductNode_POSIT1047Output_1294);

SumNode_POSIT247: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT1047Output_1294,ProductNode_POSIT943Output_1166,SumNode_POSIT247Output_1295);

ProductNode_POSIT1048: entity work.PositMult_23_6_comb_uid2(arch)
port map(v13,SumNode_POSIT247Output_1295,ProductNode_POSIT1048Output_1296);

ProductNode_POSIT1050: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1050weight,ProductNode_POSIT840Output_1039,ProductNode_POSIT1050Output_1298);

ProductNode_POSIT1087: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT258Output_1345,ProductNode_POSIT1050Output_1298,ProductNode_POSIT1087Output_1346);

ProductNode_POSIT1111: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1111weight,v14,ProductNode_POSIT1111Output_1373);

ProductNode_POSIT1112: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1112weight,vb14,ProductNode_POSIT1112Output_1374);

SumNode_POSIT262: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT1112Output_1374,ProductNode_POSIT1111Output_1373,SumNode_POSIT262Output_1375);

ProductNode_POSIT1113: entity work.PositMult_23_6_comb_uid2(arch)
port map(v15,SumNode_POSIT262Output_1375,ProductNode_POSIT1113Output_1376);

ProductNode_POSIT1114: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1114weight,ProductNode_POSIT1113Output_1376,ProductNode_POSIT1114Output_1377);

ProductNode_POSIT1115: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1115weight,v14,ProductNode_POSIT1115Output_1378);

ProductNode_POSIT1116: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1116weight,vb14,ProductNode_POSIT1116Output_1379);

SumNode_POSIT263: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT1116Output_1379,ProductNode_POSIT1115Output_1378,SumNode_POSIT263Output_1380);

ProductNode_POSIT1117: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb15,SumNode_POSIT263Output_1380,ProductNode_POSIT1117Output_1381);

ProductNode_POSIT1118: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1118weight,ProductNode_POSIT1117Output_1381,ProductNode_POSIT1118Output_1382);

SumNode_POSIT264: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT1118Output_1382,ProductNode_POSIT1114Output_1377,SumNode_POSIT264Output_1383);

ProductNode_POSIT1119: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT264Output_1383,ProductNode_POSIT901Output_1114,ProductNode_POSIT1119Output_1384);

ProductNode_POSIT1146: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1146weight,ProductNode_POSIT1113Output_1376,ProductNode_POSIT1146Output_1415);

ProductNode_POSIT1150: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1150weight,ProductNode_POSIT1117Output_1381,ProductNode_POSIT1150Output_1420);

SumNode_POSIT270: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT1150Output_1420,ProductNode_POSIT1146Output_1415,SumNode_POSIT270Output_1421);

ProductNode_POSIT1151: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT270Output_1421,ProductNode_POSIT933Output_1152,ProductNode_POSIT1151Output_1422);

SumNode_POSIT271: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT1151Output_1422,ProductNode_POSIT1119Output_1384,SumNode_POSIT271Output_1423);

ProductNode_POSIT1152: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT271Output_1423,ProductNode_POSIT1087Output_1346,ProductNode_POSIT1152Output_1424);

ProductNode_POSIT1154: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1154weight,ProductNode_POSIT944Output_1167,ProductNode_POSIT1154Output_1426);

ProductNode_POSIT1191: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT282Output_1473,ProductNode_POSIT1154Output_1426,ProductNode_POSIT1191Output_1474);

ProductNode_POSIT1218: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1218weight,ProductNode_POSIT1113Output_1376,ProductNode_POSIT1218Output_1505);

ProductNode_POSIT1222: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1222weight,ProductNode_POSIT1117Output_1381,ProductNode_POSIT1222Output_1510);

SumNode_POSIT288: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT1222Output_1510,ProductNode_POSIT1218Output_1505,SumNode_POSIT288Output_1511);

ProductNode_POSIT1223: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT288Output_1511,ProductNode_POSIT1005Output_1242,ProductNode_POSIT1223Output_1512);

ProductNode_POSIT1250: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1250weight,ProductNode_POSIT1113Output_1376,ProductNode_POSIT1250Output_1543);

ProductNode_POSIT1254: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1254weight,ProductNode_POSIT1117Output_1381,ProductNode_POSIT1254Output_1548);

SumNode_POSIT294: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT1254Output_1548,ProductNode_POSIT1250Output_1543,SumNode_POSIT294Output_1549);

ProductNode_POSIT1255: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT294Output_1549,ProductNode_POSIT1037Output_1280,ProductNode_POSIT1255Output_1550);

SumNode_POSIT295: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT1255Output_1550,ProductNode_POSIT1223Output_1512,SumNode_POSIT295Output_1551);

ProductNode_POSIT1256: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT295Output_1551,ProductNode_POSIT1191Output_1474,ProductNode_POSIT1256Output_1552);

SumNode_POSIT296: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT1256Output_1552,ProductNode_POSIT1152Output_1424,SumNode_POSIT296Output_1553);

ProductNode_POSIT1257: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb13,SumNode_POSIT296Output_1553,ProductNode_POSIT1257Output_1554);

SumNode_POSIT297: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT1257Output_1554,ProductNode_POSIT1048Output_1296,SumNode_POSIT297Output_1555);

ProductNode_POSIT1258: entity work.PositMult_23_6_comb_uid2(arch)
port map(v3,SumNode_POSIT297Output_1555,ProductNode_POSIT1258Output_1556);

ProductNode_POSIT1261: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1261weight,v2,ProductNode_POSIT1261Output_1559);

ProductNode_POSIT1278: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT302Output_1580,ProductNode_POSIT1261Output_1559,ProductNode_POSIT1278Output_1581);

ProductNode_POSIT1279: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1279weight,vb2,ProductNode_POSIT1279Output_1582);

ProductNode_POSIT1296: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT307Output_1603,ProductNode_POSIT1279Output_1582,ProductNode_POSIT1296Output_1604);

SumNode_POSIT308: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT1296Output_1604,ProductNode_POSIT1278Output_1581,SumNode_POSIT308Output_1605);

ProductNode_POSIT1297: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT308Output_1605,ProductNode_POSIT841Output_1040,ProductNode_POSIT1297Output_1606);

ProductNode_POSIT1308: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1308weight,ProductNode_POSIT468Output_579,ProductNode_POSIT1308Output_1618);

ProductNode_POSIT1318: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1318weight,ProductNode_POSIT478Output_590,ProductNode_POSIT1318Output_1629);

SumNode_POSIT311: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT1318Output_1629,ProductNode_POSIT1308Output_1618,SumNode_POSIT311Output_1630);

ProductNode_POSIT1319: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT311Output_1630,ProductNode_POSIT40Output_51,ProductNode_POSIT1319Output_1631);

ProductNode_POSIT1320: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1320weight,ProductNode_POSIT1319Output_1631,ProductNode_POSIT1320Output_1632);

ProductNode_POSIT1324: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1324weight,ProductNode_POSIT904Output_1118,ProductNode_POSIT1324Output_1637);

ProductNode_POSIT1328: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1328weight,ProductNode_POSIT908Output_1123,ProductNode_POSIT1328Output_1642);

SumNode_POSIT314: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT1328Output_1642,ProductNode_POSIT1324Output_1637,SumNode_POSIT314Output_1643);

ProductNode_POSIT1329: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT314Output_1643,ProductNode_POSIT1320Output_1632,ProductNode_POSIT1329Output_1644);

ProductNode_POSIT1340: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1340weight,ProductNode_POSIT500Output_617,ProductNode_POSIT1340Output_1656);

ProductNode_POSIT1350: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1350weight,ProductNode_POSIT510Output_628,ProductNode_POSIT1350Output_1667);

SumNode_POSIT317: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT1350Output_1667,ProductNode_POSIT1340Output_1656,SumNode_POSIT317Output_1668);

ProductNode_POSIT1351: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT317Output_1668,ProductNode_POSIT72Output_89,ProductNode_POSIT1351Output_1669);

ProductNode_POSIT1352: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1352weight,ProductNode_POSIT1351Output_1669,ProductNode_POSIT1352Output_1670);

ProductNode_POSIT1356: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1356weight,ProductNode_POSIT904Output_1118,ProductNode_POSIT1356Output_1675);

ProductNode_POSIT1360: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1360weight,ProductNode_POSIT908Output_1123,ProductNode_POSIT1360Output_1680);

SumNode_POSIT320: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT1360Output_1680,ProductNode_POSIT1356Output_1675,SumNode_POSIT320Output_1681);

ProductNode_POSIT1361: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT320Output_1681,ProductNode_POSIT1352Output_1670,ProductNode_POSIT1361Output_1682);

SumNode_POSIT321: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT1361Output_1682,ProductNode_POSIT1329Output_1644,SumNode_POSIT321Output_1683);

ProductNode_POSIT1362: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT321Output_1683,ProductNode_POSIT1297Output_1606,ProductNode_POSIT1362Output_1684);

ProductNode_POSIT1382: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT227Output_1190,ProductNode_POSIT1261Output_1559,ProductNode_POSIT1382Output_1709);

ProductNode_POSIT1400: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT232Output_1213,ProductNode_POSIT1279Output_1582,ProductNode_POSIT1400Output_1732);

SumNode_POSIT332: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT1400Output_1732,ProductNode_POSIT1382Output_1709,SumNode_POSIT332Output_1733);

ProductNode_POSIT1401: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT332Output_1733,ProductNode_POSIT945Output_1168,ProductNode_POSIT1401Output_1734);

ProductNode_POSIT1424: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1424weight,ProductNode_POSIT1319Output_1631,ProductNode_POSIT1424Output_1760);

ProductNode_POSIT1428: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1428weight,ProductNode_POSIT904Output_1118,ProductNode_POSIT1428Output_1765);

ProductNode_POSIT1432: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1432weight,ProductNode_POSIT908Output_1123,ProductNode_POSIT1432Output_1770);

SumNode_POSIT338: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT1432Output_1770,ProductNode_POSIT1428Output_1765,SumNode_POSIT338Output_1771);

ProductNode_POSIT1433: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT338Output_1771,ProductNode_POSIT1424Output_1760,ProductNode_POSIT1433Output_1772);

ProductNode_POSIT1456: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1456weight,ProductNode_POSIT1351Output_1669,ProductNode_POSIT1456Output_1798);

ProductNode_POSIT1460: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1460weight,ProductNode_POSIT904Output_1118,ProductNode_POSIT1460Output_1803);

ProductNode_POSIT1464: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1464weight,ProductNode_POSIT908Output_1123,ProductNode_POSIT1464Output_1808);

SumNode_POSIT344: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT1464Output_1808,ProductNode_POSIT1460Output_1803,SumNode_POSIT344Output_1809);

ProductNode_POSIT1465: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT344Output_1809,ProductNode_POSIT1456Output_1798,ProductNode_POSIT1465Output_1810);

SumNode_POSIT345: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT1465Output_1810,ProductNode_POSIT1433Output_1772,SumNode_POSIT345Output_1811);

ProductNode_POSIT1466: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT345Output_1811,ProductNode_POSIT1401Output_1734,ProductNode_POSIT1466Output_1812);

SumNode_POSIT346: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT1466Output_1812,ProductNode_POSIT1362Output_1684,SumNode_POSIT346Output_1813);

ProductNode_POSIT1467: entity work.PositMult_23_6_comb_uid2(arch)
port map(v13,SumNode_POSIT346Output_1813,ProductNode_POSIT1467Output_1814);

ProductNode_POSIT1506: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT357Output_1863,ProductNode_POSIT1050Output_1298,ProductNode_POSIT1506Output_1864);

ProductNode_POSIT1533: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1533weight,ProductNode_POSIT1113Output_1376,ProductNode_POSIT1533Output_1895);

ProductNode_POSIT1537: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1537weight,ProductNode_POSIT1117Output_1381,ProductNode_POSIT1537Output_1900);

SumNode_POSIT363: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT1537Output_1900,ProductNode_POSIT1533Output_1895,SumNode_POSIT363Output_1901);

ProductNode_POSIT1538: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT363Output_1901,ProductNode_POSIT1320Output_1632,ProductNode_POSIT1538Output_1902);

ProductNode_POSIT1565: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1565weight,ProductNode_POSIT1113Output_1376,ProductNode_POSIT1565Output_1933);

ProductNode_POSIT1569: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1569weight,ProductNode_POSIT1117Output_1381,ProductNode_POSIT1569Output_1938);

SumNode_POSIT369: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT1569Output_1938,ProductNode_POSIT1565Output_1933,SumNode_POSIT369Output_1939);

ProductNode_POSIT1570: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT369Output_1939,ProductNode_POSIT1352Output_1670,ProductNode_POSIT1570Output_1940);

SumNode_POSIT370: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT1570Output_1940,ProductNode_POSIT1538Output_1902,SumNode_POSIT370Output_1941);

ProductNode_POSIT1571: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT370Output_1941,ProductNode_POSIT1506Output_1864,ProductNode_POSIT1571Output_1942);

ProductNode_POSIT1610: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT381Output_1991,ProductNode_POSIT1154Output_1426,ProductNode_POSIT1610Output_1992);

ProductNode_POSIT1637: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1637weight,ProductNode_POSIT1113Output_1376,ProductNode_POSIT1637Output_2023);

ProductNode_POSIT1641: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1641weight,ProductNode_POSIT1117Output_1381,ProductNode_POSIT1641Output_2028);

SumNode_POSIT387: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT1641Output_2028,ProductNode_POSIT1637Output_2023,SumNode_POSIT387Output_2029);

ProductNode_POSIT1642: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT387Output_2029,ProductNode_POSIT1424Output_1760,ProductNode_POSIT1642Output_2030);

ProductNode_POSIT1669: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1669weight,ProductNode_POSIT1113Output_1376,ProductNode_POSIT1669Output_2061);

ProductNode_POSIT1673: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1673weight,ProductNode_POSIT1117Output_1381,ProductNode_POSIT1673Output_2066);

SumNode_POSIT393: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT1673Output_2066,ProductNode_POSIT1669Output_2061,SumNode_POSIT393Output_2067);

ProductNode_POSIT1674: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT393Output_2067,ProductNode_POSIT1456Output_1798,ProductNode_POSIT1674Output_2068);

SumNode_POSIT394: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT1674Output_2068,ProductNode_POSIT1642Output_2030,SumNode_POSIT394Output_2069);

ProductNode_POSIT1675: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT394Output_2069,ProductNode_POSIT1610Output_1992,ProductNode_POSIT1675Output_2070);

SumNode_POSIT395: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT1675Output_2070,ProductNode_POSIT1571Output_1942,SumNode_POSIT395Output_2071);

ProductNode_POSIT1676: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb13,SumNode_POSIT395Output_2071,ProductNode_POSIT1676Output_2072);

SumNode_POSIT396: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT1676Output_2072,ProductNode_POSIT1467Output_1814,SumNode_POSIT396Output_2073);

ProductNode_POSIT1677: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb3,SumNode_POSIT396Output_2073,ProductNode_POSIT1677Output_2074);

SumNode_POSIT397: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT1677Output_2074,ProductNode_POSIT1258Output_1556,SumNode_POSIT397Output_2075);

ProductNode_POSIT1678: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb4,SumNode_POSIT397Output_2075,ProductNode_POSIT1678Output_2076);

SumNode_POSIT398: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT1678Output_2076,ProductNode_POSIT839Output_1038,SumNode_POSIT398Output_2077);

ProductNode_POSIT1679: entity work.PositMult_23_6_comb_uid2(arch)
port map(v12,SumNode_POSIT398Output_2077,ProductNode_POSIT1679Output_2078);

ProductNode_POSIT1680: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1680weight,v11,ProductNode_POSIT1680Output_2079);

ProductNode_POSIT1681: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1681weight,ProductNode_POSIT1680Output_2079,ProductNode_POSIT1681Output_2080);

ProductNode_POSIT1682: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1682weight,v2,ProductNode_POSIT1682Output_2081);

ProductNode_POSIT1683: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1683weight,v7,ProductNode_POSIT1683Output_2082);

ProductNode_POSIT1684: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1684weight,vb7,ProductNode_POSIT1684Output_2083);

SumNode_POSIT399: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT1684Output_2083,ProductNode_POSIT1683Output_2082,SumNode_POSIT399Output_2084);

ProductNode_POSIT1685: entity work.PositMult_23_6_comb_uid2(arch)
port map(v1,SumNode_POSIT399Output_2084,ProductNode_POSIT1685Output_2085);

ProductNode_POSIT1686: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1686weight,v8,ProductNode_POSIT1686Output_2086);

ProductNode_POSIT1687: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1687weight,ProductNode_POSIT1686Output_2086,ProductNode_POSIT1687Output_2087);

ProductNode_POSIT1688: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1688weight,vb8,ProductNode_POSIT1688Output_2088);

ProductNode_POSIT1689: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1689weight,ProductNode_POSIT1688Output_2088,ProductNode_POSIT1689Output_2089);

SumNode_POSIT400: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT1689Output_2089,ProductNode_POSIT1687Output_2087,SumNode_POSIT400Output_2090);

ProductNode_POSIT1690: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT400Output_2090,ProductNode_POSIT1685Output_2085,ProductNode_POSIT1690Output_2091);

ProductNode_POSIT1691: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1691weight,v7,ProductNode_POSIT1691Output_2092);

ProductNode_POSIT1692: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1692weight,vb7,ProductNode_POSIT1692Output_2093);

SumNode_POSIT401: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT1692Output_2093,ProductNode_POSIT1691Output_2092,SumNode_POSIT401Output_2094);

ProductNode_POSIT1693: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb1,SumNode_POSIT401Output_2094,ProductNode_POSIT1693Output_2095);

ProductNode_POSIT1694: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1694weight,v8,ProductNode_POSIT1694Output_2096);

ProductNode_POSIT1695: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1695weight,ProductNode_POSIT1694Output_2096,ProductNode_POSIT1695Output_2097);

ProductNode_POSIT1696: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1696weight,vb8,ProductNode_POSIT1696Output_2098);

ProductNode_POSIT1697: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1697weight,ProductNode_POSIT1696Output_2098,ProductNode_POSIT1697Output_2099);

SumNode_POSIT402: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT1697Output_2099,ProductNode_POSIT1695Output_2097,SumNode_POSIT402Output_2100);

ProductNode_POSIT1698: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT402Output_2100,ProductNode_POSIT1693Output_2095,ProductNode_POSIT1698Output_2101);

SumNode_POSIT403: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT1698Output_2101,ProductNode_POSIT1690Output_2091,SumNode_POSIT403Output_2102);

ProductNode_POSIT1699: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT403Output_2102,ProductNode_POSIT1682Output_2081,ProductNode_POSIT1699Output_2103);

ProductNode_POSIT1700: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1700weight,vb2,ProductNode_POSIT1700Output_2104);

ProductNode_POSIT1704: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1704weight,v8,ProductNode_POSIT1704Output_2109);

ProductNode_POSIT1705: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1705weight,ProductNode_POSIT1704Output_2109,ProductNode_POSIT1705Output_2110);

ProductNode_POSIT1706: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1706weight,vb8,ProductNode_POSIT1706Output_2111);

ProductNode_POSIT1707: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1707weight,ProductNode_POSIT1706Output_2111,ProductNode_POSIT1707Output_2112);

SumNode_POSIT405: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT1707Output_2112,ProductNode_POSIT1705Output_2110,SumNode_POSIT405Output_2113);

ProductNode_POSIT1708: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT405Output_2113,ProductNode_POSIT1685Output_2085,ProductNode_POSIT1708Output_2114);

ProductNode_POSIT1712: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1712weight,v8,ProductNode_POSIT1712Output_2119);

ProductNode_POSIT1713: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1713weight,ProductNode_POSIT1712Output_2119,ProductNode_POSIT1713Output_2120);

ProductNode_POSIT1714: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1714weight,vb8,ProductNode_POSIT1714Output_2121);

ProductNode_POSIT1715: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1715weight,ProductNode_POSIT1714Output_2121,ProductNode_POSIT1715Output_2122);

SumNode_POSIT407: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT1715Output_2122,ProductNode_POSIT1713Output_2120,SumNode_POSIT407Output_2123);

ProductNode_POSIT1716: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT407Output_2123,ProductNode_POSIT1693Output_2095,ProductNode_POSIT1716Output_2124);

SumNode_POSIT408: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT1716Output_2124,ProductNode_POSIT1708Output_2114,SumNode_POSIT408Output_2125);

ProductNode_POSIT1717: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT408Output_2125,ProductNode_POSIT1700Output_2104,ProductNode_POSIT1717Output_2126);

SumNode_POSIT409: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT1717Output_2126,ProductNode_POSIT1699Output_2103,SumNode_POSIT409Output_2127);

ProductNode_POSIT1718: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT409Output_2127,ProductNode_POSIT1681Output_2080,ProductNode_POSIT1718Output_2128);

ProductNode_POSIT1742: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1742weight,v14,ProductNode_POSIT1742Output_2155);

ProductNode_POSIT1743: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1743weight,vb14,ProductNode_POSIT1743Output_2156);

SumNode_POSIT413: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT1743Output_2156,ProductNode_POSIT1742Output_2155,SumNode_POSIT413Output_2157);

ProductNode_POSIT1744: entity work.PositMult_23_6_comb_uid2(arch)
port map(v15,SumNode_POSIT413Output_2157,ProductNode_POSIT1744Output_2158);

ProductNode_POSIT1745: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1745weight,ProductNode_POSIT1744Output_2158,ProductNode_POSIT1745Output_2159);

ProductNode_POSIT1749: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1749weight,ProductNode_POSIT278Output_343,ProductNode_POSIT1749Output_2164);

SumNode_POSIT415: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT1749Output_2164,ProductNode_POSIT1745Output_2159,SumNode_POSIT415Output_2165);

ProductNode_POSIT1750: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT415Output_2165,ProductNode_POSIT62Output_76,ProductNode_POSIT1750Output_2166);

ProductNode_POSIT1777: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1777weight,ProductNode_POSIT1744Output_2158,ProductNode_POSIT1777Output_2197);

ProductNode_POSIT1781: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1781weight,ProductNode_POSIT278Output_343,ProductNode_POSIT1781Output_2202);

SumNode_POSIT421: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT1781Output_2202,ProductNode_POSIT1777Output_2197,SumNode_POSIT421Output_2203);

ProductNode_POSIT1782: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT421Output_2203,ProductNode_POSIT94Output_114,ProductNode_POSIT1782Output_2204);

SumNode_POSIT422: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT1782Output_2204,ProductNode_POSIT1750Output_2166,SumNode_POSIT422Output_2205);

ProductNode_POSIT1783: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT422Output_2205,ProductNode_POSIT1718Output_2128,ProductNode_POSIT1783Output_2206);

ProductNode_POSIT1784: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1784weight,vb11,ProductNode_POSIT1784Output_2207);

ProductNode_POSIT1785: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1785weight,ProductNode_POSIT1784Output_2207,ProductNode_POSIT1785Output_2208);

ProductNode_POSIT1791: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1791weight,ProductNode_POSIT1686Output_2086,ProductNode_POSIT1791Output_2215);

ProductNode_POSIT1793: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1793weight,ProductNode_POSIT1688Output_2088,ProductNode_POSIT1793Output_2217);

SumNode_POSIT424: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT1793Output_2217,ProductNode_POSIT1791Output_2215,SumNode_POSIT424Output_2218);

ProductNode_POSIT1794: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT424Output_2218,ProductNode_POSIT1685Output_2085,ProductNode_POSIT1794Output_2219);

ProductNode_POSIT1799: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1799weight,ProductNode_POSIT1694Output_2096,ProductNode_POSIT1799Output_2225);

ProductNode_POSIT1801: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1801weight,ProductNode_POSIT1696Output_2098,ProductNode_POSIT1801Output_2227);

SumNode_POSIT426: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT1801Output_2227,ProductNode_POSIT1799Output_2225,SumNode_POSIT426Output_2228);

ProductNode_POSIT1802: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT426Output_2228,ProductNode_POSIT1693Output_2095,ProductNode_POSIT1802Output_2229);

SumNode_POSIT427: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT1802Output_2229,ProductNode_POSIT1794Output_2219,SumNode_POSIT427Output_2230);

ProductNode_POSIT1803: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT427Output_2230,ProductNode_POSIT1682Output_2081,ProductNode_POSIT1803Output_2231);

ProductNode_POSIT1809: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1809weight,ProductNode_POSIT1704Output_2109,ProductNode_POSIT1809Output_2238);

ProductNode_POSIT1811: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1811weight,ProductNode_POSIT1706Output_2111,ProductNode_POSIT1811Output_2240);

SumNode_POSIT429: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT1811Output_2240,ProductNode_POSIT1809Output_2238,SumNode_POSIT429Output_2241);

ProductNode_POSIT1812: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT429Output_2241,ProductNode_POSIT1685Output_2085,ProductNode_POSIT1812Output_2242);

ProductNode_POSIT1817: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1817weight,ProductNode_POSIT1712Output_2119,ProductNode_POSIT1817Output_2248);

ProductNode_POSIT1819: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1819weight,ProductNode_POSIT1714Output_2121,ProductNode_POSIT1819Output_2250);

SumNode_POSIT431: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT1819Output_2250,ProductNode_POSIT1817Output_2248,SumNode_POSIT431Output_2251);

ProductNode_POSIT1820: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT431Output_2251,ProductNode_POSIT1693Output_2095,ProductNode_POSIT1820Output_2252);

SumNode_POSIT432: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT1820Output_2252,ProductNode_POSIT1812Output_2242,SumNode_POSIT432Output_2253);

ProductNode_POSIT1821: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT432Output_2253,ProductNode_POSIT1700Output_2104,ProductNode_POSIT1821Output_2254);

SumNode_POSIT433: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT1821Output_2254,ProductNode_POSIT1803Output_2231,SumNode_POSIT433Output_2255);

ProductNode_POSIT1822: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT433Output_2255,ProductNode_POSIT1785Output_2208,ProductNode_POSIT1822Output_2256);

ProductNode_POSIT1849: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1849weight,ProductNode_POSIT1744Output_2158,ProductNode_POSIT1849Output_2287);

ProductNode_POSIT1853: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1853weight,ProductNode_POSIT278Output_343,ProductNode_POSIT1853Output_2292);

SumNode_POSIT439: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT1853Output_2292,ProductNode_POSIT1849Output_2287,SumNode_POSIT439Output_2293);

ProductNode_POSIT1854: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT439Output_2293,ProductNode_POSIT166Output_204,ProductNode_POSIT1854Output_2294);

ProductNode_POSIT1881: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1881weight,ProductNode_POSIT1744Output_2158,ProductNode_POSIT1881Output_2325);

ProductNode_POSIT1885: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1885weight,ProductNode_POSIT278Output_343,ProductNode_POSIT1885Output_2330);

SumNode_POSIT445: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT1885Output_2330,ProductNode_POSIT1881Output_2325,SumNode_POSIT445Output_2331);

ProductNode_POSIT1886: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT445Output_2331,ProductNode_POSIT198Output_242,ProductNode_POSIT1886Output_2332);

SumNode_POSIT446: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT1886Output_2332,ProductNode_POSIT1854Output_2294,SumNode_POSIT446Output_2333);

ProductNode_POSIT1887: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT446Output_2333,ProductNode_POSIT1822Output_2256,ProductNode_POSIT1887Output_2334);

SumNode_POSIT447: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT1887Output_2334,ProductNode_POSIT1783Output_2206,SumNode_POSIT447Output_2335);

ProductNode_POSIT1888: entity work.PositMult_23_6_comb_uid2(arch)
port map(v13,SumNode_POSIT447Output_2335,ProductNode_POSIT1888Output_2336);

ProductNode_POSIT1890: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1890weight,ProductNode_POSIT1680Output_2079,ProductNode_POSIT1890Output_2338);

ProductNode_POSIT1927: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT458Output_2385,ProductNode_POSIT1890Output_2338,ProductNode_POSIT1927Output_2386);

ProductNode_POSIT1951: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1951weight,v14,ProductNode_POSIT1951Output_2413);

ProductNode_POSIT1952: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1952weight,vb14,ProductNode_POSIT1952Output_2414);

SumNode_POSIT462: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT1952Output_2414,ProductNode_POSIT1951Output_2413,SumNode_POSIT462Output_2415);

ProductNode_POSIT1953: entity work.PositMult_23_6_comb_uid2(arch)
port map(v15,SumNode_POSIT462Output_2415,ProductNode_POSIT1953Output_2416);

ProductNode_POSIT1954: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1954weight,ProductNode_POSIT1953Output_2416,ProductNode_POSIT1954Output_2417);

ProductNode_POSIT1955: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1955weight,v14,ProductNode_POSIT1955Output_2418);

ProductNode_POSIT1956: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1956weight,vb14,ProductNode_POSIT1956Output_2419);

SumNode_POSIT463: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT1956Output_2419,ProductNode_POSIT1955Output_2418,SumNode_POSIT463Output_2420);

ProductNode_POSIT1957: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb15,SumNode_POSIT463Output_2420,ProductNode_POSIT1957Output_2421);

ProductNode_POSIT1958: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1958weight,ProductNode_POSIT1957Output_2421,ProductNode_POSIT1958Output_2422);

SumNode_POSIT464: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT1958Output_2422,ProductNode_POSIT1954Output_2417,SumNode_POSIT464Output_2423);

ProductNode_POSIT1959: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT464Output_2423,ProductNode_POSIT62Output_76,ProductNode_POSIT1959Output_2424);

ProductNode_POSIT1986: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1986weight,ProductNode_POSIT1953Output_2416,ProductNode_POSIT1986Output_2455);

ProductNode_POSIT1990: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1990weight,ProductNode_POSIT1957Output_2421,ProductNode_POSIT1990Output_2460);

SumNode_POSIT470: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT1990Output_2460,ProductNode_POSIT1986Output_2455,SumNode_POSIT470Output_2461);

ProductNode_POSIT1991: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT470Output_2461,ProductNode_POSIT94Output_114,ProductNode_POSIT1991Output_2462);

SumNode_POSIT471: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT1991Output_2462,ProductNode_POSIT1959Output_2424,SumNode_POSIT471Output_2463);

ProductNode_POSIT1992: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT471Output_2463,ProductNode_POSIT1927Output_2386,ProductNode_POSIT1992Output_2464);

ProductNode_POSIT1994: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT1994weight,ProductNode_POSIT1784Output_2207,ProductNode_POSIT1994Output_2466);

ProductNode_POSIT2031: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT482Output_2513,ProductNode_POSIT1994Output_2466,ProductNode_POSIT2031Output_2514);

ProductNode_POSIT2058: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT2058weight,ProductNode_POSIT1953Output_2416,ProductNode_POSIT2058Output_2545);

ProductNode_POSIT2062: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT2062weight,ProductNode_POSIT1957Output_2421,ProductNode_POSIT2062Output_2550);

SumNode_POSIT488: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT2062Output_2550,ProductNode_POSIT2058Output_2545,SumNode_POSIT488Output_2551);

ProductNode_POSIT2063: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT488Output_2551,ProductNode_POSIT166Output_204,ProductNode_POSIT2063Output_2552);

ProductNode_POSIT2090: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT2090weight,ProductNode_POSIT1953Output_2416,ProductNode_POSIT2090Output_2583);

ProductNode_POSIT2094: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT2094weight,ProductNode_POSIT1957Output_2421,ProductNode_POSIT2094Output_2588);

SumNode_POSIT494: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT2094Output_2588,ProductNode_POSIT2090Output_2583,SumNode_POSIT494Output_2589);

ProductNode_POSIT2095: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT494Output_2589,ProductNode_POSIT198Output_242,ProductNode_POSIT2095Output_2590);

SumNode_POSIT495: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT2095Output_2590,ProductNode_POSIT2063Output_2552,SumNode_POSIT495Output_2591);

ProductNode_POSIT2096: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT495Output_2591,ProductNode_POSIT2031Output_2514,ProductNode_POSIT2096Output_2592);

SumNode_POSIT496: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT2096Output_2592,ProductNode_POSIT1992Output_2464,SumNode_POSIT496Output_2593);

ProductNode_POSIT2097: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb13,SumNode_POSIT496Output_2593,ProductNode_POSIT2097Output_2594);

SumNode_POSIT497: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT2097Output_2594,ProductNode_POSIT1888Output_2336,SumNode_POSIT497Output_2595);

ProductNode_POSIT2098: entity work.PositMult_23_6_comb_uid2(arch)
port map(v3,SumNode_POSIT497Output_2595,ProductNode_POSIT2098Output_2596);

ProductNode_POSIT2101: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT2101weight,v2,ProductNode_POSIT2101Output_2599);

ProductNode_POSIT2118: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT502Output_2620,ProductNode_POSIT2101Output_2599,ProductNode_POSIT2118Output_2621);

ProductNode_POSIT2119: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT2119weight,vb2,ProductNode_POSIT2119Output_2622);

ProductNode_POSIT2136: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT507Output_2643,ProductNode_POSIT2119Output_2622,ProductNode_POSIT2136Output_2644);

SumNode_POSIT508: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT2136Output_2644,ProductNode_POSIT2118Output_2621,SumNode_POSIT508Output_2645);

ProductNode_POSIT2137: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT508Output_2645,ProductNode_POSIT1681Output_2080,ProductNode_POSIT2137Output_2646);

ProductNode_POSIT2164: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT2164weight,ProductNode_POSIT1744Output_2158,ProductNode_POSIT2164Output_2677);

ProductNode_POSIT2168: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT2168weight,ProductNode_POSIT278Output_343,ProductNode_POSIT2168Output_2682);

SumNode_POSIT514: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT2168Output_2682,ProductNode_POSIT2164Output_2677,SumNode_POSIT514Output_2683);

ProductNode_POSIT2169: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT514Output_2683,ProductNode_POSIT481Output_594,ProductNode_POSIT2169Output_2684);

ProductNode_POSIT2196: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT2196weight,ProductNode_POSIT1744Output_2158,ProductNode_POSIT2196Output_2715);

ProductNode_POSIT2200: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT2200weight,ProductNode_POSIT278Output_343,ProductNode_POSIT2200Output_2720);

SumNode_POSIT520: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT2200Output_2720,ProductNode_POSIT2196Output_2715,SumNode_POSIT520Output_2721);

ProductNode_POSIT2201: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT520Output_2721,ProductNode_POSIT513Output_632,ProductNode_POSIT2201Output_2722);

SumNode_POSIT521: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT2201Output_2722,ProductNode_POSIT2169Output_2684,SumNode_POSIT521Output_2723);

ProductNode_POSIT2202: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT521Output_2723,ProductNode_POSIT2137Output_2646,ProductNode_POSIT2202Output_2724);

ProductNode_POSIT2222: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT427Output_2230,ProductNode_POSIT2101Output_2599,ProductNode_POSIT2222Output_2749);

ProductNode_POSIT2240: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT432Output_2253,ProductNode_POSIT2119Output_2622,ProductNode_POSIT2240Output_2772);

SumNode_POSIT532: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT2240Output_2772,ProductNode_POSIT2222Output_2749,SumNode_POSIT532Output_2773);

ProductNode_POSIT2241: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT532Output_2773,ProductNode_POSIT1785Output_2208,ProductNode_POSIT2241Output_2774);

ProductNode_POSIT2268: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT2268weight,ProductNode_POSIT1744Output_2158,ProductNode_POSIT2268Output_2805);

ProductNode_POSIT2272: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT2272weight,ProductNode_POSIT278Output_343,ProductNode_POSIT2272Output_2810);

SumNode_POSIT538: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT2272Output_2810,ProductNode_POSIT2268Output_2805,SumNode_POSIT538Output_2811);

ProductNode_POSIT2273: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT538Output_2811,ProductNode_POSIT585Output_722,ProductNode_POSIT2273Output_2812);

ProductNode_POSIT2300: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT2300weight,ProductNode_POSIT1744Output_2158,ProductNode_POSIT2300Output_2843);

ProductNode_POSIT2304: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT2304weight,ProductNode_POSIT278Output_343,ProductNode_POSIT2304Output_2848);

SumNode_POSIT544: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT2304Output_2848,ProductNode_POSIT2300Output_2843,SumNode_POSIT544Output_2849);

ProductNode_POSIT2305: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT544Output_2849,ProductNode_POSIT617Output_760,ProductNode_POSIT2305Output_2850);

SumNode_POSIT545: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT2305Output_2850,ProductNode_POSIT2273Output_2812,SumNode_POSIT545Output_2851);

ProductNode_POSIT2306: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT545Output_2851,ProductNode_POSIT2241Output_2774,ProductNode_POSIT2306Output_2852);

SumNode_POSIT546: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT2306Output_2852,ProductNode_POSIT2202Output_2724,SumNode_POSIT546Output_2853);

ProductNode_POSIT2307: entity work.PositMult_23_6_comb_uid2(arch)
port map(v13,SumNode_POSIT546Output_2853,ProductNode_POSIT2307Output_2854);

ProductNode_POSIT2346: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT557Output_2903,ProductNode_POSIT1890Output_2338,ProductNode_POSIT2346Output_2904);

ProductNode_POSIT2373: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT2373weight,ProductNode_POSIT1953Output_2416,ProductNode_POSIT2373Output_2935);

ProductNode_POSIT2377: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT2377weight,ProductNode_POSIT1957Output_2421,ProductNode_POSIT2377Output_2940);

SumNode_POSIT563: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT2377Output_2940,ProductNode_POSIT2373Output_2935,SumNode_POSIT563Output_2941);

ProductNode_POSIT2378: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT563Output_2941,ProductNode_POSIT481Output_594,ProductNode_POSIT2378Output_2942);

ProductNode_POSIT2405: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT2405weight,ProductNode_POSIT1953Output_2416,ProductNode_POSIT2405Output_2973);

ProductNode_POSIT2409: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT2409weight,ProductNode_POSIT1957Output_2421,ProductNode_POSIT2409Output_2978);

SumNode_POSIT569: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT2409Output_2978,ProductNode_POSIT2405Output_2973,SumNode_POSIT569Output_2979);

ProductNode_POSIT2410: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT569Output_2979,ProductNode_POSIT513Output_632,ProductNode_POSIT2410Output_2980);

SumNode_POSIT570: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT2410Output_2980,ProductNode_POSIT2378Output_2942,SumNode_POSIT570Output_2981);

ProductNode_POSIT2411: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT570Output_2981,ProductNode_POSIT2346Output_2904,ProductNode_POSIT2411Output_2982);

ProductNode_POSIT2450: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT581Output_3031,ProductNode_POSIT1994Output_2466,ProductNode_POSIT2450Output_3032);

ProductNode_POSIT2477: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT2477weight,ProductNode_POSIT1953Output_2416,ProductNode_POSIT2477Output_3063);

ProductNode_POSIT2481: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT2481weight,ProductNode_POSIT1957Output_2421,ProductNode_POSIT2481Output_3068);

SumNode_POSIT587: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT2481Output_3068,ProductNode_POSIT2477Output_3063,SumNode_POSIT587Output_3069);

ProductNode_POSIT2482: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT587Output_3069,ProductNode_POSIT585Output_722,ProductNode_POSIT2482Output_3070);

ProductNode_POSIT2509: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT2509weight,ProductNode_POSIT1953Output_2416,ProductNode_POSIT2509Output_3101);

ProductNode_POSIT2513: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT2513weight,ProductNode_POSIT1957Output_2421,ProductNode_POSIT2513Output_3106);

SumNode_POSIT593: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT2513Output_3106,ProductNode_POSIT2509Output_3101,SumNode_POSIT593Output_3107);

ProductNode_POSIT2514: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT593Output_3107,ProductNode_POSIT617Output_760,ProductNode_POSIT2514Output_3108);

SumNode_POSIT594: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT2514Output_3108,ProductNode_POSIT2482Output_3070,SumNode_POSIT594Output_3109);

ProductNode_POSIT2515: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT594Output_3109,ProductNode_POSIT2450Output_3032,ProductNode_POSIT2515Output_3110);

SumNode_POSIT595: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT2515Output_3110,ProductNode_POSIT2411Output_2982,SumNode_POSIT595Output_3111);

ProductNode_POSIT2516: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb13,SumNode_POSIT595Output_3111,ProductNode_POSIT2516Output_3112);

SumNode_POSIT596: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT2516Output_3112,ProductNode_POSIT2307Output_2854,SumNode_POSIT596Output_3113);

ProductNode_POSIT2517: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb3,SumNode_POSIT596Output_3113,ProductNode_POSIT2517Output_3114);

SumNode_POSIT597: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT2517Output_3114,ProductNode_POSIT2098Output_2596,SumNode_POSIT597Output_3115);

ProductNode_POSIT2518: entity work.PositMult_23_6_comb_uid2(arch)
port map(v4,SumNode_POSIT597Output_3115,ProductNode_POSIT2518Output_3116);

ProductNode_POSIT2519: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT2519weight,v11,ProductNode_POSIT2519Output_3117);

ProductNode_POSIT2520: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT2520weight,ProductNode_POSIT2519Output_3117,ProductNode_POSIT2520Output_3118);

ProductNode_POSIT2521: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT2521weight,v2,ProductNode_POSIT2521Output_3119);

ProductNode_POSIT2522: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT2522weight,v7,ProductNode_POSIT2522Output_3120);

ProductNode_POSIT2523: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT2523weight,vb7,ProductNode_POSIT2523Output_3121);

SumNode_POSIT598: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT2523Output_3121,ProductNode_POSIT2522Output_3120,SumNode_POSIT598Output_3122);

ProductNode_POSIT2524: entity work.PositMult_23_6_comb_uid2(arch)
port map(v1,SumNode_POSIT598Output_3122,ProductNode_POSIT2524Output_3123);

ProductNode_POSIT2529: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT599Output_3128,ProductNode_POSIT2524Output_3123,ProductNode_POSIT2529Output_3129);

ProductNode_POSIT2530: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT2530weight,v7,ProductNode_POSIT2530Output_3130);

ProductNode_POSIT2531: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT2531weight,vb7,ProductNode_POSIT2531Output_3131);

SumNode_POSIT600: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT2531Output_3131,ProductNode_POSIT2530Output_3130,SumNode_POSIT600Output_3132);

ProductNode_POSIT2532: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb1,SumNode_POSIT600Output_3132,ProductNode_POSIT2532Output_3133);

ProductNode_POSIT2537: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT601Output_3138,ProductNode_POSIT2532Output_3133,ProductNode_POSIT2537Output_3139);

SumNode_POSIT602: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT2537Output_3139,ProductNode_POSIT2529Output_3129,SumNode_POSIT602Output_3140);

ProductNode_POSIT2538: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT602Output_3140,ProductNode_POSIT2521Output_3119,ProductNode_POSIT2538Output_3141);

ProductNode_POSIT2539: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT2539weight,vb2,ProductNode_POSIT2539Output_3142);

ProductNode_POSIT2547: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT405Output_2113,ProductNode_POSIT2524Output_3123,ProductNode_POSIT2547Output_3152);

ProductNode_POSIT2555: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT407Output_2123,ProductNode_POSIT2532Output_3133,ProductNode_POSIT2555Output_3162);

SumNode_POSIT607: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT2555Output_3162,ProductNode_POSIT2547Output_3152,SumNode_POSIT607Output_3163);

ProductNode_POSIT2556: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT607Output_3163,ProductNode_POSIT2539Output_3142,ProductNode_POSIT2556Output_3164);

SumNode_POSIT608: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT2556Output_3164,ProductNode_POSIT2538Output_3141,SumNode_POSIT608Output_3165);

ProductNode_POSIT2557: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT608Output_3165,ProductNode_POSIT2520Output_3118,ProductNode_POSIT2557Output_3166);

ProductNode_POSIT2581: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT2581weight,v14,ProductNode_POSIT2581Output_3193);

ProductNode_POSIT2582: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT2582weight,vb14,ProductNode_POSIT2582Output_3194);

SumNode_POSIT612: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT2582Output_3194,ProductNode_POSIT2581Output_3193,SumNode_POSIT612Output_3195);

ProductNode_POSIT2583: entity work.PositMult_23_6_comb_uid2(arch)
port map(v15,SumNode_POSIT612Output_3195,ProductNode_POSIT2583Output_3196);

ProductNode_POSIT2584: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT2584weight,ProductNode_POSIT2583Output_3196,ProductNode_POSIT2584Output_3197);

ProductNode_POSIT2585: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT2585weight,v14,ProductNode_POSIT2585Output_3198);

ProductNode_POSIT2586: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT2586weight,vb14,ProductNode_POSIT2586Output_3199);

SumNode_POSIT613: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT2586Output_3199,ProductNode_POSIT2585Output_3198,SumNode_POSIT613Output_3200);

ProductNode_POSIT2587: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb15,SumNode_POSIT613Output_3200,ProductNode_POSIT2587Output_3201);

ProductNode_POSIT2588: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT2588weight,ProductNode_POSIT2587Output_3201,ProductNode_POSIT2588Output_3202);

SumNode_POSIT614: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT2588Output_3202,ProductNode_POSIT2584Output_3197,SumNode_POSIT614Output_3203);

ProductNode_POSIT2589: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT614Output_3203,ProductNode_POSIT901Output_1114,ProductNode_POSIT2589Output_3204);

ProductNode_POSIT2616: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT2616weight,ProductNode_POSIT2583Output_3196,ProductNode_POSIT2616Output_3235);

ProductNode_POSIT2620: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT2620weight,ProductNode_POSIT2587Output_3201,ProductNode_POSIT2620Output_3240);

SumNode_POSIT620: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT2620Output_3240,ProductNode_POSIT2616Output_3235,SumNode_POSIT620Output_3241);

ProductNode_POSIT2621: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT620Output_3241,ProductNode_POSIT933Output_1152,ProductNode_POSIT2621Output_3242);

SumNode_POSIT621: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT2621Output_3242,ProductNode_POSIT2589Output_3204,SumNode_POSIT621Output_3243);

ProductNode_POSIT2622: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT621Output_3243,ProductNode_POSIT2557Output_3166,ProductNode_POSIT2622Output_3244);

ProductNode_POSIT2623: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT2623weight,vb11,ProductNode_POSIT2623Output_3245);

ProductNode_POSIT2624: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT2624weight,ProductNode_POSIT2623Output_3245,ProductNode_POSIT2624Output_3246);

ProductNode_POSIT2633: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT424Output_2218,ProductNode_POSIT2524Output_3123,ProductNode_POSIT2633Output_3257);

ProductNode_POSIT2641: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT426Output_2228,ProductNode_POSIT2532Output_3133,ProductNode_POSIT2641Output_3267);

SumNode_POSIT626: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT2641Output_3267,ProductNode_POSIT2633Output_3257,SumNode_POSIT626Output_3268);

ProductNode_POSIT2642: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT626Output_3268,ProductNode_POSIT2521Output_3119,ProductNode_POSIT2642Output_3269);

ProductNode_POSIT2651: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT429Output_2241,ProductNode_POSIT2524Output_3123,ProductNode_POSIT2651Output_3280);

ProductNode_POSIT2659: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT431Output_2251,ProductNode_POSIT2532Output_3133,ProductNode_POSIT2659Output_3290);

SumNode_POSIT631: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT2659Output_3290,ProductNode_POSIT2651Output_3280,SumNode_POSIT631Output_3291);

ProductNode_POSIT2660: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT631Output_3291,ProductNode_POSIT2539Output_3142,ProductNode_POSIT2660Output_3292);

SumNode_POSIT632: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT2660Output_3292,ProductNode_POSIT2642Output_3269,SumNode_POSIT632Output_3293);

ProductNode_POSIT2661: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT632Output_3293,ProductNode_POSIT2624Output_3246,ProductNode_POSIT2661Output_3294);

ProductNode_POSIT2688: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT2688weight,ProductNode_POSIT2583Output_3196,ProductNode_POSIT2688Output_3325);

ProductNode_POSIT2692: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT2692weight,ProductNode_POSIT2587Output_3201,ProductNode_POSIT2692Output_3330);

SumNode_POSIT638: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT2692Output_3330,ProductNode_POSIT2688Output_3325,SumNode_POSIT638Output_3331);

ProductNode_POSIT2693: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT638Output_3331,ProductNode_POSIT1005Output_1242,ProductNode_POSIT2693Output_3332);

ProductNode_POSIT2720: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT2720weight,ProductNode_POSIT2583Output_3196,ProductNode_POSIT2720Output_3363);

ProductNode_POSIT2724: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT2724weight,ProductNode_POSIT2587Output_3201,ProductNode_POSIT2724Output_3368);

SumNode_POSIT644: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT2724Output_3368,ProductNode_POSIT2720Output_3363,SumNode_POSIT644Output_3369);

ProductNode_POSIT2725: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT644Output_3369,ProductNode_POSIT1037Output_1280,ProductNode_POSIT2725Output_3370);

SumNode_POSIT645: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT2725Output_3370,ProductNode_POSIT2693Output_3332,SumNode_POSIT645Output_3371);

ProductNode_POSIT2726: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT645Output_3371,ProductNode_POSIT2661Output_3294,ProductNode_POSIT2726Output_3372);

SumNode_POSIT646: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT2726Output_3372,ProductNode_POSIT2622Output_3244,SumNode_POSIT646Output_3373);

ProductNode_POSIT2727: entity work.PositMult_23_6_comb_uid2(arch)
port map(v13,SumNode_POSIT646Output_3373,ProductNode_POSIT2727Output_3374);

ProductNode_POSIT2729: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT2729weight,ProductNode_POSIT2519Output_3117,ProductNode_POSIT2729Output_3376);

ProductNode_POSIT2766: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT657Output_3423,ProductNode_POSIT2729Output_3376,ProductNode_POSIT2766Output_3424);

ProductNode_POSIT2790: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT2790weight,v14,ProductNode_POSIT2790Output_3451);

ProductNode_POSIT2791: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT2791weight,vb14,ProductNode_POSIT2791Output_3452);

SumNode_POSIT661: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT2791Output_3452,ProductNode_POSIT2790Output_3451,SumNode_POSIT661Output_3453);

ProductNode_POSIT2792: entity work.PositMult_23_6_comb_uid2(arch)
port map(v15,SumNode_POSIT661Output_3453,ProductNode_POSIT2792Output_3454);

ProductNode_POSIT2793: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT2793weight,ProductNode_POSIT2792Output_3454,ProductNode_POSIT2793Output_3455);

ProductNode_POSIT2794: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT2794weight,v14,ProductNode_POSIT2794Output_3456);

ProductNode_POSIT2795: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT2795weight,vb14,ProductNode_POSIT2795Output_3457);

SumNode_POSIT662: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT2795Output_3457,ProductNode_POSIT2794Output_3456,SumNode_POSIT662Output_3458);

ProductNode_POSIT2796: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb15,SumNode_POSIT662Output_3458,ProductNode_POSIT2796Output_3459);

ProductNode_POSIT2797: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT2797weight,ProductNode_POSIT2796Output_3459,ProductNode_POSIT2797Output_3460);

SumNode_POSIT663: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT2797Output_3460,ProductNode_POSIT2793Output_3455,SumNode_POSIT663Output_3461);

ProductNode_POSIT2798: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT663Output_3461,ProductNode_POSIT901Output_1114,ProductNode_POSIT2798Output_3462);

ProductNode_POSIT2825: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT2825weight,ProductNode_POSIT2792Output_3454,ProductNode_POSIT2825Output_3493);

ProductNode_POSIT2829: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT2829weight,ProductNode_POSIT2796Output_3459,ProductNode_POSIT2829Output_3498);

SumNode_POSIT669: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT2829Output_3498,ProductNode_POSIT2825Output_3493,SumNode_POSIT669Output_3499);

ProductNode_POSIT2830: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT669Output_3499,ProductNode_POSIT933Output_1152,ProductNode_POSIT2830Output_3500);

SumNode_POSIT670: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT2830Output_3500,ProductNode_POSIT2798Output_3462,SumNode_POSIT670Output_3501);

ProductNode_POSIT2831: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT670Output_3501,ProductNode_POSIT2766Output_3424,ProductNode_POSIT2831Output_3502);

ProductNode_POSIT2833: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT2833weight,ProductNode_POSIT2623Output_3245,ProductNode_POSIT2833Output_3504);

ProductNode_POSIT2870: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT681Output_3551,ProductNode_POSIT2833Output_3504,ProductNode_POSIT2870Output_3552);

ProductNode_POSIT2897: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT2897weight,ProductNode_POSIT2792Output_3454,ProductNode_POSIT2897Output_3583);

ProductNode_POSIT2901: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT2901weight,ProductNode_POSIT2796Output_3459,ProductNode_POSIT2901Output_3588);

SumNode_POSIT687: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT2901Output_3588,ProductNode_POSIT2897Output_3583,SumNode_POSIT687Output_3589);

ProductNode_POSIT2902: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT687Output_3589,ProductNode_POSIT1005Output_1242,ProductNode_POSIT2902Output_3590);

ProductNode_POSIT2929: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT2929weight,ProductNode_POSIT2792Output_3454,ProductNode_POSIT2929Output_3621);

ProductNode_POSIT2933: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT2933weight,ProductNode_POSIT2796Output_3459,ProductNode_POSIT2933Output_3626);

SumNode_POSIT693: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT2933Output_3626,ProductNode_POSIT2929Output_3621,SumNode_POSIT693Output_3627);

ProductNode_POSIT2934: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT693Output_3627,ProductNode_POSIT1037Output_1280,ProductNode_POSIT2934Output_3628);

SumNode_POSIT694: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT2934Output_3628,ProductNode_POSIT2902Output_3590,SumNode_POSIT694Output_3629);

ProductNode_POSIT2935: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT694Output_3629,ProductNode_POSIT2870Output_3552,ProductNode_POSIT2935Output_3630);

SumNode_POSIT695: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT2935Output_3630,ProductNode_POSIT2831Output_3502,SumNode_POSIT695Output_3631);

ProductNode_POSIT2936: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb13,SumNode_POSIT695Output_3631,ProductNode_POSIT2936Output_3632);

SumNode_POSIT696: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT2936Output_3632,ProductNode_POSIT2727Output_3374,SumNode_POSIT696Output_3633);

ProductNode_POSIT2937: entity work.PositMult_23_6_comb_uid2(arch)
port map(v3,SumNode_POSIT696Output_3633,ProductNode_POSIT2937Output_3634);

ProductNode_POSIT2940: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT2940weight,v2,ProductNode_POSIT2940Output_3637);

ProductNode_POSIT2957: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT701Output_3658,ProductNode_POSIT2940Output_3637,ProductNode_POSIT2957Output_3659);

ProductNode_POSIT2958: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT2958weight,vb2,ProductNode_POSIT2958Output_3660);

ProductNode_POSIT2975: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT706Output_3681,ProductNode_POSIT2958Output_3660,ProductNode_POSIT2975Output_3682);

SumNode_POSIT707: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT2975Output_3682,ProductNode_POSIT2957Output_3659,SumNode_POSIT707Output_3683);

ProductNode_POSIT2976: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT707Output_3683,ProductNode_POSIT2520Output_3118,ProductNode_POSIT2976Output_3684);

ProductNode_POSIT3003: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT3003weight,ProductNode_POSIT2583Output_3196,ProductNode_POSIT3003Output_3715);

ProductNode_POSIT3007: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT3007weight,ProductNode_POSIT2587Output_3201,ProductNode_POSIT3007Output_3720);

SumNode_POSIT713: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT3007Output_3720,ProductNode_POSIT3003Output_3715,SumNode_POSIT713Output_3721);

ProductNode_POSIT3008: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT713Output_3721,ProductNode_POSIT1320Output_1632,ProductNode_POSIT3008Output_3722);

ProductNode_POSIT3035: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT3035weight,ProductNode_POSIT2583Output_3196,ProductNode_POSIT3035Output_3753);

ProductNode_POSIT3039: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT3039weight,ProductNode_POSIT2587Output_3201,ProductNode_POSIT3039Output_3758);

SumNode_POSIT719: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT3039Output_3758,ProductNode_POSIT3035Output_3753,SumNode_POSIT719Output_3759);

ProductNode_POSIT3040: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT719Output_3759,ProductNode_POSIT1352Output_1670,ProductNode_POSIT3040Output_3760);

SumNode_POSIT720: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT3040Output_3760,ProductNode_POSIT3008Output_3722,SumNode_POSIT720Output_3761);

ProductNode_POSIT3041: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT720Output_3761,ProductNode_POSIT2976Output_3684,ProductNode_POSIT3041Output_3762);

ProductNode_POSIT3061: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT626Output_3268,ProductNode_POSIT2940Output_3637,ProductNode_POSIT3061Output_3787);

ProductNode_POSIT3079: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT631Output_3291,ProductNode_POSIT2958Output_3660,ProductNode_POSIT3079Output_3810);

SumNode_POSIT731: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT3079Output_3810,ProductNode_POSIT3061Output_3787,SumNode_POSIT731Output_3811);

ProductNode_POSIT3080: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT731Output_3811,ProductNode_POSIT2624Output_3246,ProductNode_POSIT3080Output_3812);

ProductNode_POSIT3107: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT3107weight,ProductNode_POSIT2583Output_3196,ProductNode_POSIT3107Output_3843);

ProductNode_POSIT3111: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT3111weight,ProductNode_POSIT2587Output_3201,ProductNode_POSIT3111Output_3848);

SumNode_POSIT737: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT3111Output_3848,ProductNode_POSIT3107Output_3843,SumNode_POSIT737Output_3849);

ProductNode_POSIT3112: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT737Output_3849,ProductNode_POSIT1424Output_1760,ProductNode_POSIT3112Output_3850);

ProductNode_POSIT3139: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT3139weight,ProductNode_POSIT2583Output_3196,ProductNode_POSIT3139Output_3881);

ProductNode_POSIT3143: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT3143weight,ProductNode_POSIT2587Output_3201,ProductNode_POSIT3143Output_3886);

SumNode_POSIT743: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT3143Output_3886,ProductNode_POSIT3139Output_3881,SumNode_POSIT743Output_3887);

ProductNode_POSIT3144: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT743Output_3887,ProductNode_POSIT1456Output_1798,ProductNode_POSIT3144Output_3888);

SumNode_POSIT744: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT3144Output_3888,ProductNode_POSIT3112Output_3850,SumNode_POSIT744Output_3889);

ProductNode_POSIT3145: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT744Output_3889,ProductNode_POSIT3080Output_3812,ProductNode_POSIT3145Output_3890);

SumNode_POSIT745: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT3145Output_3890,ProductNode_POSIT3041Output_3762,SumNode_POSIT745Output_3891);

ProductNode_POSIT3146: entity work.PositMult_23_6_comb_uid2(arch)
port map(v13,SumNode_POSIT745Output_3891,ProductNode_POSIT3146Output_3892);

ProductNode_POSIT3185: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT756Output_3941,ProductNode_POSIT2729Output_3376,ProductNode_POSIT3185Output_3942);

ProductNode_POSIT3212: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT3212weight,ProductNode_POSIT2792Output_3454,ProductNode_POSIT3212Output_3973);

ProductNode_POSIT3216: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT3216weight,ProductNode_POSIT2796Output_3459,ProductNode_POSIT3216Output_3978);

SumNode_POSIT762: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT3216Output_3978,ProductNode_POSIT3212Output_3973,SumNode_POSIT762Output_3979);

ProductNode_POSIT3217: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT762Output_3979,ProductNode_POSIT1320Output_1632,ProductNode_POSIT3217Output_3980);

ProductNode_POSIT3244: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT3244weight,ProductNode_POSIT2792Output_3454,ProductNode_POSIT3244Output_4011);

ProductNode_POSIT3248: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT3248weight,ProductNode_POSIT2796Output_3459,ProductNode_POSIT3248Output_4016);

SumNode_POSIT768: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT3248Output_4016,ProductNode_POSIT3244Output_4011,SumNode_POSIT768Output_4017);

ProductNode_POSIT3249: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT768Output_4017,ProductNode_POSIT1352Output_1670,ProductNode_POSIT3249Output_4018);

SumNode_POSIT769: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT3249Output_4018,ProductNode_POSIT3217Output_3980,SumNode_POSIT769Output_4019);

ProductNode_POSIT3250: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT769Output_4019,ProductNode_POSIT3185Output_3942,ProductNode_POSIT3250Output_4020);

ProductNode_POSIT3289: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT780Output_4069,ProductNode_POSIT2833Output_3504,ProductNode_POSIT3289Output_4070);

ProductNode_POSIT3316: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT3316weight,ProductNode_POSIT2792Output_3454,ProductNode_POSIT3316Output_4101);

ProductNode_POSIT3320: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT3320weight,ProductNode_POSIT2796Output_3459,ProductNode_POSIT3320Output_4106);

SumNode_POSIT786: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT3320Output_4106,ProductNode_POSIT3316Output_4101,SumNode_POSIT786Output_4107);

ProductNode_POSIT3321: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT786Output_4107,ProductNode_POSIT1424Output_1760,ProductNode_POSIT3321Output_4108);

ProductNode_POSIT3348: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT3348weight,ProductNode_POSIT2792Output_3454,ProductNode_POSIT3348Output_4139);

ProductNode_POSIT3352: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT3352weight,ProductNode_POSIT2796Output_3459,ProductNode_POSIT3352Output_4144);

SumNode_POSIT792: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT3352Output_4144,ProductNode_POSIT3348Output_4139,SumNode_POSIT792Output_4145);

ProductNode_POSIT3353: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT792Output_4145,ProductNode_POSIT1456Output_1798,ProductNode_POSIT3353Output_4146);

SumNode_POSIT793: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT3353Output_4146,ProductNode_POSIT3321Output_4108,SumNode_POSIT793Output_4147);

ProductNode_POSIT3354: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT793Output_4147,ProductNode_POSIT3289Output_4070,ProductNode_POSIT3354Output_4148);

SumNode_POSIT794: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT3354Output_4148,ProductNode_POSIT3250Output_4020,SumNode_POSIT794Output_4149);

ProductNode_POSIT3355: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb13,SumNode_POSIT794Output_4149,ProductNode_POSIT3355Output_4150);

SumNode_POSIT795: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT3355Output_4150,ProductNode_POSIT3146Output_3892,SumNode_POSIT795Output_4151);

ProductNode_POSIT3356: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb3,SumNode_POSIT795Output_4151,ProductNode_POSIT3356Output_4152);

SumNode_POSIT796: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT3356Output_4152,ProductNode_POSIT2937Output_3634,SumNode_POSIT796Output_4153);

ProductNode_POSIT3357: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb4,SumNode_POSIT796Output_4153,ProductNode_POSIT3357Output_4154);

SumNode_POSIT797: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT3357Output_4154,ProductNode_POSIT2518Output_3116,SumNode_POSIT797Output_4155);

ProductNode_POSIT3358: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb12,SumNode_POSIT797Output_4155,ProductNode_POSIT3358Output_4156);

SumNode_POSIT798: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT3358Output_4156,ProductNode_POSIT1679Output_2078,SumNode_POSIT798Output_4157);

ProductNode_POSIT3359: entity work.PositMult_23_6_comb_uid2(arch)
port map(v6,SumNode_POSIT798Output_4157,ProductNode_POSIT3359Output_4158);

ProductNode_POSIT3361: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT3361weight,ProductNode_POSIT1Output_1,ProductNode_POSIT3361Output_4160);

ProductNode_POSIT3363: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT3363weight,v7,ProductNode_POSIT3363Output_4162);

ProductNode_POSIT3364: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT3364weight,vb7,ProductNode_POSIT3364Output_4163);

SumNode_POSIT799: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT3364Output_4163,ProductNode_POSIT3363Output_4162,SumNode_POSIT799Output_4164);

ProductNode_POSIT3365: entity work.PositMult_23_6_comb_uid2(arch)
port map(v1,SumNode_POSIT799Output_4164,ProductNode_POSIT3365Output_4165);

ProductNode_POSIT3370: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT800Output_4170,ProductNode_POSIT3365Output_4165,ProductNode_POSIT3370Output_4171);

ProductNode_POSIT3371: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT3371weight,v7,ProductNode_POSIT3371Output_4172);

ProductNode_POSIT3372: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT3372weight,vb7,ProductNode_POSIT3372Output_4173);

SumNode_POSIT801: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT3372Output_4173,ProductNode_POSIT3371Output_4172,SumNode_POSIT801Output_4174);

ProductNode_POSIT3373: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb1,SumNode_POSIT801Output_4174,ProductNode_POSIT3373Output_4175);

ProductNode_POSIT3378: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT802Output_4180,ProductNode_POSIT3373Output_4175,ProductNode_POSIT3378Output_4181);

SumNode_POSIT803: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT3378Output_4181,ProductNode_POSIT3370Output_4171,SumNode_POSIT803Output_4182);

ProductNode_POSIT3379: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT803Output_4182,ProductNode_POSIT3Output_3,ProductNode_POSIT3379Output_4183);

ProductNode_POSIT3388: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT6Output_35,ProductNode_POSIT3365Output_4165,ProductNode_POSIT3388Output_4194);

ProductNode_POSIT3396: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT8Output_45,ProductNode_POSIT3373Output_4175,ProductNode_POSIT3396Output_4204);

SumNode_POSIT808: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT3396Output_4204,ProductNode_POSIT3388Output_4194,SumNode_POSIT808Output_4205);

ProductNode_POSIT3397: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT808Output_4205,ProductNode_POSIT21Output_26,ProductNode_POSIT3397Output_4206);

SumNode_POSIT809: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT3397Output_4206,ProductNode_POSIT3379Output_4183,SumNode_POSIT809Output_4207);

ProductNode_POSIT3398: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT809Output_4207,ProductNode_POSIT3361Output_4160,ProductNode_POSIT3398Output_4208);

ProductNode_POSIT3401: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT3401weight,ProductNode_POSIT41Output_52,ProductNode_POSIT3401Output_4211);

ProductNode_POSIT3402: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT3402weight,ProductNode_POSIT3401Output_4211,ProductNode_POSIT3402Output_4212);

ProductNode_POSIT3403: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT3403weight,ProductNode_POSIT3402Output_4212,ProductNode_POSIT3403Output_4213);

ProductNode_POSIT3405: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT3405weight,ProductNode_POSIT45Output_56,ProductNode_POSIT3405Output_4215);

ProductNode_POSIT3406: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT3406weight,ProductNode_POSIT3405Output_4215,ProductNode_POSIT3406Output_4216);

ProductNode_POSIT3407: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT3407weight,ProductNode_POSIT3406Output_4216,ProductNode_POSIT3407Output_4217);

SumNode_POSIT810: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT3407Output_4217,ProductNode_POSIT3403Output_4213,SumNode_POSIT810Output_4218);

ProductNode_POSIT3408: entity work.PositMult_23_6_comb_uid2(arch)
port map(v16,SumNode_POSIT810Output_4218,ProductNode_POSIT3408Output_4219);

ProductNode_POSIT3409: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT3409weight,ProductNode_POSIT3408Output_4219,ProductNode_POSIT3409Output_4220);

ProductNode_POSIT3412: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT3412weight,ProductNode_POSIT3401Output_4211,ProductNode_POSIT3412Output_4223);

ProductNode_POSIT3413: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT3413weight,ProductNode_POSIT3412Output_4223,ProductNode_POSIT3413Output_4224);

ProductNode_POSIT3416: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT3416weight,ProductNode_POSIT3405Output_4215,ProductNode_POSIT3416Output_4227);

ProductNode_POSIT3417: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT3417weight,ProductNode_POSIT3416Output_4227,ProductNode_POSIT3417Output_4228);

SumNode_POSIT811: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT3417Output_4228,ProductNode_POSIT3413Output_4224,SumNode_POSIT811Output_4229);

ProductNode_POSIT3418: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb16,SumNode_POSIT811Output_4229,ProductNode_POSIT3418Output_4230);

ProductNode_POSIT3419: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT3419weight,ProductNode_POSIT3418Output_4230,ProductNode_POSIT3419Output_4231);

SumNode_POSIT812: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT3419Output_4231,ProductNode_POSIT3409Output_4220,SumNode_POSIT812Output_4232);

ProductNode_POSIT3420: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT812Output_4232,ProductNode_POSIT40Output_51,ProductNode_POSIT3420Output_4233);

ProductNode_POSIT3421: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT3421weight,ProductNode_POSIT3420Output_4233,ProductNode_POSIT3421Output_4234);

ProductNode_POSIT3430: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT815Output_4245,ProductNode_POSIT3421Output_4234,ProductNode_POSIT3430Output_4246);

ProductNode_POSIT3433: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT3433weight,ProductNode_POSIT73Output_90,ProductNode_POSIT3433Output_4249);

ProductNode_POSIT3434: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT3434weight,ProductNode_POSIT3433Output_4249,ProductNode_POSIT3434Output_4250);

ProductNode_POSIT3435: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT3435weight,ProductNode_POSIT3434Output_4250,ProductNode_POSIT3435Output_4251);

ProductNode_POSIT3437: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT3437weight,ProductNode_POSIT77Output_94,ProductNode_POSIT3437Output_4253);

ProductNode_POSIT3438: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT3438weight,ProductNode_POSIT3437Output_4253,ProductNode_POSIT3438Output_4254);

ProductNode_POSIT3439: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT3439weight,ProductNode_POSIT3438Output_4254,ProductNode_POSIT3439Output_4255);

SumNode_POSIT816: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT3439Output_4255,ProductNode_POSIT3435Output_4251,SumNode_POSIT816Output_4256);

ProductNode_POSIT3440: entity work.PositMult_23_6_comb_uid2(arch)
port map(v16,SumNode_POSIT816Output_4256,ProductNode_POSIT3440Output_4257);

ProductNode_POSIT3441: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT3441weight,ProductNode_POSIT3440Output_4257,ProductNode_POSIT3441Output_4258);

ProductNode_POSIT3444: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT3444weight,ProductNode_POSIT3433Output_4249,ProductNode_POSIT3444Output_4261);

ProductNode_POSIT3445: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT3445weight,ProductNode_POSIT3444Output_4261,ProductNode_POSIT3445Output_4262);

ProductNode_POSIT3448: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT3448weight,ProductNode_POSIT3437Output_4253,ProductNode_POSIT3448Output_4265);

ProductNode_POSIT3449: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT3449weight,ProductNode_POSIT3448Output_4265,ProductNode_POSIT3449Output_4266);

SumNode_POSIT817: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT3449Output_4266,ProductNode_POSIT3445Output_4262,SumNode_POSIT817Output_4267);

ProductNode_POSIT3450: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb16,SumNode_POSIT817Output_4267,ProductNode_POSIT3450Output_4268);

ProductNode_POSIT3451: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT3451weight,ProductNode_POSIT3450Output_4268,ProductNode_POSIT3451Output_4269);

SumNode_POSIT818: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT3451Output_4269,ProductNode_POSIT3441Output_4258,SumNode_POSIT818Output_4270);

ProductNode_POSIT3452: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT818Output_4270,ProductNode_POSIT72Output_89,ProductNode_POSIT3452Output_4271);

ProductNode_POSIT3453: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT3453weight,ProductNode_POSIT3452Output_4271,ProductNode_POSIT3453Output_4272);

ProductNode_POSIT3462: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT821Output_4283,ProductNode_POSIT3453Output_4272,ProductNode_POSIT3462Output_4284);

SumNode_POSIT822: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT3462Output_4284,ProductNode_POSIT3430Output_4246,SumNode_POSIT822Output_4285);

ProductNode_POSIT3463: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT822Output_4285,ProductNode_POSIT3398Output_4208,ProductNode_POSIT3463Output_4286);

ProductNode_POSIT3465: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT3465weight,ProductNode_POSIT105Output_129,ProductNode_POSIT3465Output_4288);

ProductNode_POSIT3474: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT25Output_140,ProductNode_POSIT3365Output_4165,ProductNode_POSIT3474Output_4299);

ProductNode_POSIT3482: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT27Output_150,ProductNode_POSIT3373Output_4175,ProductNode_POSIT3482Output_4309);

SumNode_POSIT827: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT3482Output_4309,ProductNode_POSIT3474Output_4299,SumNode_POSIT827Output_4310);

ProductNode_POSIT3483: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT827Output_4310,ProductNode_POSIT3Output_3,ProductNode_POSIT3483Output_4311);

ProductNode_POSIT3492: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT30Output_163,ProductNode_POSIT3365Output_4165,ProductNode_POSIT3492Output_4322);

ProductNode_POSIT3500: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT32Output_173,ProductNode_POSIT3373Output_4175,ProductNode_POSIT3500Output_4332);

SumNode_POSIT832: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT3500Output_4332,ProductNode_POSIT3492Output_4322,SumNode_POSIT832Output_4333);

ProductNode_POSIT3501: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT832Output_4333,ProductNode_POSIT21Output_26,ProductNode_POSIT3501Output_4334);

SumNode_POSIT833: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT3501Output_4334,ProductNode_POSIT3483Output_4311,SumNode_POSIT833Output_4335);

ProductNode_POSIT3502: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT833Output_4335,ProductNode_POSIT3465Output_4288,ProductNode_POSIT3502Output_4336);

ProductNode_POSIT3525: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT3525weight,ProductNode_POSIT3420Output_4233,ProductNode_POSIT3525Output_4362);

ProductNode_POSIT3534: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT839Output_4373,ProductNode_POSIT3525Output_4362,ProductNode_POSIT3534Output_4374);

ProductNode_POSIT3557: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT3557weight,ProductNode_POSIT3452Output_4271,ProductNode_POSIT3557Output_4400);

ProductNode_POSIT3566: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT845Output_4411,ProductNode_POSIT3557Output_4400,ProductNode_POSIT3566Output_4412);

SumNode_POSIT846: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT3566Output_4412,ProductNode_POSIT3534Output_4374,SumNode_POSIT846Output_4413);

ProductNode_POSIT3567: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT846Output_4413,ProductNode_POSIT3502Output_4336,ProductNode_POSIT3567Output_4414);

SumNode_POSIT847: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT3567Output_4414,ProductNode_POSIT3463Output_4286,SumNode_POSIT847Output_4415);

ProductNode_POSIT3568: entity work.PositMult_23_6_comb_uid2(arch)
port map(v13,SumNode_POSIT847Output_4415,ProductNode_POSIT3568Output_4416);

ProductNode_POSIT3570: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT3570weight,ProductNode_POSIT1Output_1,ProductNode_POSIT3570Output_4418);

ProductNode_POSIT3607: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT858Output_4465,ProductNode_POSIT3570Output_4418,ProductNode_POSIT3607Output_4466);

ProductNode_POSIT3639: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT65Output_345,ProductNode_POSIT3421Output_4234,ProductNode_POSIT3639Output_4504);

ProductNode_POSIT3671: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT71Output_383,ProductNode_POSIT3453Output_4272,ProductNode_POSIT3671Output_4542);

SumNode_POSIT871: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT3671Output_4542,ProductNode_POSIT3639Output_4504,SumNode_POSIT871Output_4543);

ProductNode_POSIT3672: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT871Output_4543,ProductNode_POSIT3607Output_4466,ProductNode_POSIT3672Output_4544);

ProductNode_POSIT3674: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT3674weight,ProductNode_POSIT105Output_129,ProductNode_POSIT3674Output_4546);

ProductNode_POSIT3711: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT882Output_4593,ProductNode_POSIT3674Output_4546,ProductNode_POSIT3711Output_4594);

ProductNode_POSIT3743: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT89Output_473,ProductNode_POSIT3525Output_4362,ProductNode_POSIT3743Output_4632);

ProductNode_POSIT3775: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT95Output_511,ProductNode_POSIT3557Output_4400,ProductNode_POSIT3775Output_4670);

SumNode_POSIT895: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT3775Output_4670,ProductNode_POSIT3743Output_4632,SumNode_POSIT895Output_4671);

ProductNode_POSIT3776: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT895Output_4671,ProductNode_POSIT3711Output_4594,ProductNode_POSIT3776Output_4672);

SumNode_POSIT896: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT3776Output_4672,ProductNode_POSIT3672Output_4544,SumNode_POSIT896Output_4673);

ProductNode_POSIT3777: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb13,SumNode_POSIT896Output_4673,ProductNode_POSIT3777Output_4674);

SumNode_POSIT897: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT3777Output_4674,ProductNode_POSIT3568Output_4416,SumNode_POSIT897Output_4675);

ProductNode_POSIT3778: entity work.PositMult_23_6_comb_uid2(arch)
port map(v3,SumNode_POSIT897Output_4675,ProductNode_POSIT3778Output_4676);

ProductNode_POSIT3798: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT902Output_4700,ProductNode_POSIT422Output_521,ProductNode_POSIT3798Output_4701);

ProductNode_POSIT3816: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT907Output_4723,ProductNode_POSIT440Output_544,ProductNode_POSIT3816Output_4724);

SumNode_POSIT908: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT3816Output_4724,ProductNode_POSIT3798Output_4701,SumNode_POSIT908Output_4725);

ProductNode_POSIT3817: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT908Output_4725,ProductNode_POSIT3361Output_4160,ProductNode_POSIT3817Output_4726);

ProductNode_POSIT3822: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT3822weight,ProductNode_POSIT3402Output_4212,ProductNode_POSIT3822Output_4731);

ProductNode_POSIT3826: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT3826weight,ProductNode_POSIT3406Output_4216,ProductNode_POSIT3826Output_4735);

SumNode_POSIT909: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT3826Output_4735,ProductNode_POSIT3822Output_4731,SumNode_POSIT909Output_4736);

ProductNode_POSIT3827: entity work.PositMult_23_6_comb_uid2(arch)
port map(v16,SumNode_POSIT909Output_4736,ProductNode_POSIT3827Output_4737);

ProductNode_POSIT3828: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT3828weight,ProductNode_POSIT3827Output_4737,ProductNode_POSIT3828Output_4738);

ProductNode_POSIT3832: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT3832weight,ProductNode_POSIT3412Output_4223,ProductNode_POSIT3832Output_4742);

ProductNode_POSIT3836: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT3836weight,ProductNode_POSIT3416Output_4227,ProductNode_POSIT3836Output_4746);

SumNode_POSIT910: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT3836Output_4746,ProductNode_POSIT3832Output_4742,SumNode_POSIT910Output_4747);

ProductNode_POSIT3837: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb16,SumNode_POSIT910Output_4747,ProductNode_POSIT3837Output_4748);

ProductNode_POSIT3838: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT3838weight,ProductNode_POSIT3837Output_4748,ProductNode_POSIT3838Output_4749);

SumNode_POSIT911: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT3838Output_4749,ProductNode_POSIT3828Output_4738,SumNode_POSIT911Output_4750);

ProductNode_POSIT3839: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT911Output_4750,ProductNode_POSIT40Output_51,ProductNode_POSIT3839Output_4751);

ProductNode_POSIT3840: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT3840weight,ProductNode_POSIT3839Output_4751,ProductNode_POSIT3840Output_4752);

ProductNode_POSIT3849: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT914Output_4763,ProductNode_POSIT3840Output_4752,ProductNode_POSIT3849Output_4764);

ProductNode_POSIT3854: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT3854weight,ProductNode_POSIT3434Output_4250,ProductNode_POSIT3854Output_4769);

ProductNode_POSIT3858: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT3858weight,ProductNode_POSIT3438Output_4254,ProductNode_POSIT3858Output_4773);

SumNode_POSIT915: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT3858Output_4773,ProductNode_POSIT3854Output_4769,SumNode_POSIT915Output_4774);

ProductNode_POSIT3859: entity work.PositMult_23_6_comb_uid2(arch)
port map(v16,SumNode_POSIT915Output_4774,ProductNode_POSIT3859Output_4775);

ProductNode_POSIT3860: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT3860weight,ProductNode_POSIT3859Output_4775,ProductNode_POSIT3860Output_4776);

ProductNode_POSIT3864: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT3864weight,ProductNode_POSIT3444Output_4261,ProductNode_POSIT3864Output_4780);

ProductNode_POSIT3868: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT3868weight,ProductNode_POSIT3448Output_4265,ProductNode_POSIT3868Output_4784);

SumNode_POSIT916: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT3868Output_4784,ProductNode_POSIT3864Output_4780,SumNode_POSIT916Output_4785);

ProductNode_POSIT3869: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb16,SumNode_POSIT916Output_4785,ProductNode_POSIT3869Output_4786);

ProductNode_POSIT3870: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT3870weight,ProductNode_POSIT3869Output_4786,ProductNode_POSIT3870Output_4787);

SumNode_POSIT917: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT3870Output_4787,ProductNode_POSIT3860Output_4776,SumNode_POSIT917Output_4788);

ProductNode_POSIT3871: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT917Output_4788,ProductNode_POSIT72Output_89,ProductNode_POSIT3871Output_4789);

ProductNode_POSIT3872: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT3872weight,ProductNode_POSIT3871Output_4789,ProductNode_POSIT3872Output_4790);

ProductNode_POSIT3881: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT920Output_4801,ProductNode_POSIT3872Output_4790,ProductNode_POSIT3881Output_4802);

SumNode_POSIT921: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT3881Output_4802,ProductNode_POSIT3849Output_4764,SumNode_POSIT921Output_4803);

ProductNode_POSIT3882: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT921Output_4803,ProductNode_POSIT3817Output_4726,ProductNode_POSIT3882Output_4804);

ProductNode_POSIT3902: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT926Output_4828,ProductNode_POSIT422Output_521,ProductNode_POSIT3902Output_4829);

ProductNode_POSIT3920: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT931Output_4851,ProductNode_POSIT440Output_544,ProductNode_POSIT3920Output_4852);

SumNode_POSIT932: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT3920Output_4852,ProductNode_POSIT3902Output_4829,SumNode_POSIT932Output_4853);

ProductNode_POSIT3921: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT932Output_4853,ProductNode_POSIT3465Output_4288,ProductNode_POSIT3921Output_4854);

ProductNode_POSIT3944: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT3944weight,ProductNode_POSIT3839Output_4751,ProductNode_POSIT3944Output_4880);

ProductNode_POSIT3953: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT938Output_4891,ProductNode_POSIT3944Output_4880,ProductNode_POSIT3953Output_4892);

ProductNode_POSIT3976: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT3976weight,ProductNode_POSIT3871Output_4789,ProductNode_POSIT3976Output_4918);

ProductNode_POSIT3985: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT944Output_4929,ProductNode_POSIT3976Output_4918,ProductNode_POSIT3985Output_4930);

SumNode_POSIT945: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT3985Output_4930,ProductNode_POSIT3953Output_4892,SumNode_POSIT945Output_4931);

ProductNode_POSIT3986: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT945Output_4931,ProductNode_POSIT3921Output_4854,ProductNode_POSIT3986Output_4932);

SumNode_POSIT946: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT3986Output_4932,ProductNode_POSIT3882Output_4804,SumNode_POSIT946Output_4933);

ProductNode_POSIT3987: entity work.PositMult_23_6_comb_uid2(arch)
port map(v13,SumNode_POSIT946Output_4933,ProductNode_POSIT3987Output_4934);

ProductNode_POSIT4026: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT957Output_4983,ProductNode_POSIT3570Output_4418,ProductNode_POSIT4026Output_4984);

ProductNode_POSIT4058: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT164Output_863,ProductNode_POSIT3840Output_4752,ProductNode_POSIT4058Output_5022);

ProductNode_POSIT4090: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT170Output_901,ProductNode_POSIT3872Output_4790,ProductNode_POSIT4090Output_5060);

SumNode_POSIT970: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT4090Output_5060,ProductNode_POSIT4058Output_5022,SumNode_POSIT970Output_5061);

ProductNode_POSIT4091: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT970Output_5061,ProductNode_POSIT4026Output_4984,ProductNode_POSIT4091Output_5062);

ProductNode_POSIT4130: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT981Output_5111,ProductNode_POSIT3674Output_4546,ProductNode_POSIT4130Output_5112);

ProductNode_POSIT4162: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT188Output_991,ProductNode_POSIT3944Output_4880,ProductNode_POSIT4162Output_5150);

ProductNode_POSIT4194: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT194Output_1029,ProductNode_POSIT3976Output_4918,ProductNode_POSIT4194Output_5188);

SumNode_POSIT994: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT4194Output_5188,ProductNode_POSIT4162Output_5150,SumNode_POSIT994Output_5189);

ProductNode_POSIT4195: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT994Output_5189,ProductNode_POSIT4130Output_5112,ProductNode_POSIT4195Output_5190);

SumNode_POSIT995: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT4195Output_5190,ProductNode_POSIT4091Output_5062,SumNode_POSIT995Output_5191);

ProductNode_POSIT4196: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb13,SumNode_POSIT995Output_5191,ProductNode_POSIT4196Output_5192);

SumNode_POSIT996: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT4196Output_5192,ProductNode_POSIT3987Output_4934,SumNode_POSIT996Output_5193);

ProductNode_POSIT4197: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb3,SumNode_POSIT996Output_5193,ProductNode_POSIT4197Output_5194);

SumNode_POSIT997: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT4197Output_5194,ProductNode_POSIT3778Output_4676,SumNode_POSIT997Output_5195);

ProductNode_POSIT4198: entity work.PositMult_23_6_comb_uid2(arch)
port map(v4,SumNode_POSIT997Output_5195,ProductNode_POSIT4198Output_5196);

ProductNode_POSIT4200: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT4200weight,ProductNode_POSIT840Output_1039,ProductNode_POSIT4200Output_5198);

ProductNode_POSIT4202: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT4202weight,v7,ProductNode_POSIT4202Output_5200);

ProductNode_POSIT4203: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT4203weight,vb7,ProductNode_POSIT4203Output_5201);

SumNode_POSIT998: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT4203Output_5201,ProductNode_POSIT4202Output_5200,SumNode_POSIT998Output_5202);

ProductNode_POSIT4204: entity work.PositMult_23_6_comb_uid2(arch)
port map(v1,SumNode_POSIT998Output_5202,ProductNode_POSIT4204Output_5203);

ProductNode_POSIT4209: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT999Output_5208,ProductNode_POSIT4204Output_5203,ProductNode_POSIT4209Output_5209);

ProductNode_POSIT4210: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT4210weight,v7,ProductNode_POSIT4210Output_5210);

ProductNode_POSIT4211: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT4211weight,vb7,ProductNode_POSIT4211Output_5211);

SumNode_POSIT1000: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT4211Output_5211,ProductNode_POSIT4210Output_5210,SumNode_POSIT1000Output_5212);

ProductNode_POSIT4212: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb1,SumNode_POSIT1000Output_5212,ProductNode_POSIT4212Output_5213);

ProductNode_POSIT4217: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1001Output_5218,ProductNode_POSIT4212Output_5213,ProductNode_POSIT4217Output_5219);

SumNode_POSIT1002: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT4217Output_5219,ProductNode_POSIT4209Output_5209,SumNode_POSIT1002Output_5220);

ProductNode_POSIT4218: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1002Output_5220,ProductNode_POSIT842Output_1041,ProductNode_POSIT4218Output_5221);

ProductNode_POSIT4227: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT6Output_35,ProductNode_POSIT4204Output_5203,ProductNode_POSIT4227Output_5232);

ProductNode_POSIT4235: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT8Output_45,ProductNode_POSIT4212Output_5213,ProductNode_POSIT4235Output_5242);

SumNode_POSIT1007: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT4235Output_5242,ProductNode_POSIT4227Output_5232,SumNode_POSIT1007Output_5243);

ProductNode_POSIT4236: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1007Output_5243,ProductNode_POSIT860Output_1064,ProductNode_POSIT4236Output_5244);

SumNode_POSIT1008: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT4236Output_5244,ProductNode_POSIT4218Output_5221,SumNode_POSIT1008Output_5245);

ProductNode_POSIT4237: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1008Output_5245,ProductNode_POSIT4200Output_5198,ProductNode_POSIT4237Output_5246);

ProductNode_POSIT4248: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT4248weight,ProductNode_POSIT3408Output_4219,ProductNode_POSIT4248Output_5258);

ProductNode_POSIT4258: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT4258weight,ProductNode_POSIT3418Output_4230,ProductNode_POSIT4258Output_5269);

SumNode_POSIT1011: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT4258Output_5269,ProductNode_POSIT4248Output_5258,SumNode_POSIT1011Output_5270);

ProductNode_POSIT4259: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1011Output_5270,ProductNode_POSIT40Output_51,ProductNode_POSIT4259Output_5271);

ProductNode_POSIT4260: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT4260weight,ProductNode_POSIT4259Output_5271,ProductNode_POSIT4260Output_5272);

ProductNode_POSIT4269: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1014Output_5283,ProductNode_POSIT4260Output_5272,ProductNode_POSIT4269Output_5284);

ProductNode_POSIT4280: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT4280weight,ProductNode_POSIT3440Output_4257,ProductNode_POSIT4280Output_5296);

ProductNode_POSIT4290: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT4290weight,ProductNode_POSIT3450Output_4268,ProductNode_POSIT4290Output_5307);

SumNode_POSIT1017: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT4290Output_5307,ProductNode_POSIT4280Output_5296,SumNode_POSIT1017Output_5308);

ProductNode_POSIT4291: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1017Output_5308,ProductNode_POSIT72Output_89,ProductNode_POSIT4291Output_5309);

ProductNode_POSIT4292: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT4292weight,ProductNode_POSIT4291Output_5309,ProductNode_POSIT4292Output_5310);

ProductNode_POSIT4301: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1020Output_5321,ProductNode_POSIT4292Output_5310,ProductNode_POSIT4301Output_5322);

SumNode_POSIT1021: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT4301Output_5322,ProductNode_POSIT4269Output_5284,SumNode_POSIT1021Output_5323);

ProductNode_POSIT4302: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1021Output_5323,ProductNode_POSIT4237Output_5246,ProductNode_POSIT4302Output_5324);

ProductNode_POSIT4304: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT4304weight,ProductNode_POSIT944Output_1167,ProductNode_POSIT4304Output_5326);

ProductNode_POSIT4313: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT25Output_140,ProductNode_POSIT4204Output_5203,ProductNode_POSIT4313Output_5337);

ProductNode_POSIT4321: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT27Output_150,ProductNode_POSIT4212Output_5213,ProductNode_POSIT4321Output_5347);

SumNode_POSIT1026: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT4321Output_5347,ProductNode_POSIT4313Output_5337,SumNode_POSIT1026Output_5348);

ProductNode_POSIT4322: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1026Output_5348,ProductNode_POSIT842Output_1041,ProductNode_POSIT4322Output_5349);

ProductNode_POSIT4331: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT30Output_163,ProductNode_POSIT4204Output_5203,ProductNode_POSIT4331Output_5360);

ProductNode_POSIT4339: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT32Output_173,ProductNode_POSIT4212Output_5213,ProductNode_POSIT4339Output_5370);

SumNode_POSIT1031: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT4339Output_5370,ProductNode_POSIT4331Output_5360,SumNode_POSIT1031Output_5371);

ProductNode_POSIT4340: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1031Output_5371,ProductNode_POSIT860Output_1064,ProductNode_POSIT4340Output_5372);

SumNode_POSIT1032: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT4340Output_5372,ProductNode_POSIT4322Output_5349,SumNode_POSIT1032Output_5373);

ProductNode_POSIT4341: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1032Output_5373,ProductNode_POSIT4304Output_5326,ProductNode_POSIT4341Output_5374);

ProductNode_POSIT4364: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT4364weight,ProductNode_POSIT4259Output_5271,ProductNode_POSIT4364Output_5400);

ProductNode_POSIT4373: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1038Output_5411,ProductNode_POSIT4364Output_5400,ProductNode_POSIT4373Output_5412);

ProductNode_POSIT4396: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT4396weight,ProductNode_POSIT4291Output_5309,ProductNode_POSIT4396Output_5438);

ProductNode_POSIT4405: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1044Output_5449,ProductNode_POSIT4396Output_5438,ProductNode_POSIT4405Output_5450);

SumNode_POSIT1045: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT4405Output_5450,ProductNode_POSIT4373Output_5412,SumNode_POSIT1045Output_5451);

ProductNode_POSIT4406: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1045Output_5451,ProductNode_POSIT4341Output_5374,ProductNode_POSIT4406Output_5452);

SumNode_POSIT1046: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT4406Output_5452,ProductNode_POSIT4302Output_5324,SumNode_POSIT1046Output_5453);

ProductNode_POSIT4407: entity work.PositMult_23_6_comb_uid2(arch)
port map(v13,SumNode_POSIT1046Output_5453,ProductNode_POSIT4407Output_5454);

ProductNode_POSIT4409: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT4409weight,ProductNode_POSIT840Output_1039,ProductNode_POSIT4409Output_5456);

ProductNode_POSIT4446: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1057Output_5503,ProductNode_POSIT4409Output_5456,ProductNode_POSIT4446Output_5504);

ProductNode_POSIT4478: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT264Output_1383,ProductNode_POSIT4260Output_5272,ProductNode_POSIT4478Output_5542);

ProductNode_POSIT4510: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT270Output_1421,ProductNode_POSIT4292Output_5310,ProductNode_POSIT4510Output_5580);

SumNode_POSIT1070: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT4510Output_5580,ProductNode_POSIT4478Output_5542,SumNode_POSIT1070Output_5581);

ProductNode_POSIT4511: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1070Output_5581,ProductNode_POSIT4446Output_5504,ProductNode_POSIT4511Output_5582);

ProductNode_POSIT4513: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT4513weight,ProductNode_POSIT944Output_1167,ProductNode_POSIT4513Output_5584);

ProductNode_POSIT4550: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1081Output_5631,ProductNode_POSIT4513Output_5584,ProductNode_POSIT4550Output_5632);

ProductNode_POSIT4582: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT288Output_1511,ProductNode_POSIT4364Output_5400,ProductNode_POSIT4582Output_5670);

ProductNode_POSIT4614: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT294Output_1549,ProductNode_POSIT4396Output_5438,ProductNode_POSIT4614Output_5708);

SumNode_POSIT1094: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT4614Output_5708,ProductNode_POSIT4582Output_5670,SumNode_POSIT1094Output_5709);

ProductNode_POSIT4615: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1094Output_5709,ProductNode_POSIT4550Output_5632,ProductNode_POSIT4615Output_5710);

SumNode_POSIT1095: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT4615Output_5710,ProductNode_POSIT4511Output_5582,SumNode_POSIT1095Output_5711);

ProductNode_POSIT4616: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb13,SumNode_POSIT1095Output_5711,ProductNode_POSIT4616Output_5712);

SumNode_POSIT1096: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT4616Output_5712,ProductNode_POSIT4407Output_5454,SumNode_POSIT1096Output_5713);

ProductNode_POSIT4617: entity work.PositMult_23_6_comb_uid2(arch)
port map(v3,SumNode_POSIT1096Output_5713,ProductNode_POSIT4617Output_5714);

ProductNode_POSIT4637: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1101Output_5738,ProductNode_POSIT1261Output_1559,ProductNode_POSIT4637Output_5739);

ProductNode_POSIT4655: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1106Output_5761,ProductNode_POSIT1279Output_1582,ProductNode_POSIT4655Output_5762);

SumNode_POSIT1107: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT4655Output_5762,ProductNode_POSIT4637Output_5739,SumNode_POSIT1107Output_5763);

ProductNode_POSIT4656: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1107Output_5763,ProductNode_POSIT4200Output_5198,ProductNode_POSIT4656Output_5764);

ProductNode_POSIT4667: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT4667weight,ProductNode_POSIT3827Output_4737,ProductNode_POSIT4667Output_5776);

ProductNode_POSIT4677: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT4677weight,ProductNode_POSIT3837Output_4748,ProductNode_POSIT4677Output_5787);

SumNode_POSIT1110: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT4677Output_5787,ProductNode_POSIT4667Output_5776,SumNode_POSIT1110Output_5788);

ProductNode_POSIT4678: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1110Output_5788,ProductNode_POSIT40Output_51,ProductNode_POSIT4678Output_5789);

ProductNode_POSIT4679: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT4679weight,ProductNode_POSIT4678Output_5789,ProductNode_POSIT4679Output_5790);

ProductNode_POSIT4688: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1113Output_5801,ProductNode_POSIT4679Output_5790,ProductNode_POSIT4688Output_5802);

ProductNode_POSIT4699: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT4699weight,ProductNode_POSIT3859Output_4775,ProductNode_POSIT4699Output_5814);

ProductNode_POSIT4709: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT4709weight,ProductNode_POSIT3869Output_4786,ProductNode_POSIT4709Output_5825);

SumNode_POSIT1116: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT4709Output_5825,ProductNode_POSIT4699Output_5814,SumNode_POSIT1116Output_5826);

ProductNode_POSIT4710: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1116Output_5826,ProductNode_POSIT72Output_89,ProductNode_POSIT4710Output_5827);

ProductNode_POSIT4711: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT4711weight,ProductNode_POSIT4710Output_5827,ProductNode_POSIT4711Output_5828);

ProductNode_POSIT4720: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1119Output_5839,ProductNode_POSIT4711Output_5828,ProductNode_POSIT4720Output_5840);

SumNode_POSIT1120: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT4720Output_5840,ProductNode_POSIT4688Output_5802,SumNode_POSIT1120Output_5841);

ProductNode_POSIT4721: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1120Output_5841,ProductNode_POSIT4656Output_5764,ProductNode_POSIT4721Output_5842);

ProductNode_POSIT4741: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1125Output_5866,ProductNode_POSIT1261Output_1559,ProductNode_POSIT4741Output_5867);

ProductNode_POSIT4759: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1130Output_5889,ProductNode_POSIT1279Output_1582,ProductNode_POSIT4759Output_5890);

SumNode_POSIT1131: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT4759Output_5890,ProductNode_POSIT4741Output_5867,SumNode_POSIT1131Output_5891);

ProductNode_POSIT4760: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1131Output_5891,ProductNode_POSIT4304Output_5326,ProductNode_POSIT4760Output_5892);

ProductNode_POSIT4783: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT4783weight,ProductNode_POSIT4678Output_5789,ProductNode_POSIT4783Output_5918);

ProductNode_POSIT4792: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1137Output_5929,ProductNode_POSIT4783Output_5918,ProductNode_POSIT4792Output_5930);

ProductNode_POSIT4815: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT4815weight,ProductNode_POSIT4710Output_5827,ProductNode_POSIT4815Output_5956);

ProductNode_POSIT4824: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1143Output_5967,ProductNode_POSIT4815Output_5956,ProductNode_POSIT4824Output_5968);

SumNode_POSIT1144: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT4824Output_5968,ProductNode_POSIT4792Output_5930,SumNode_POSIT1144Output_5969);

ProductNode_POSIT4825: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1144Output_5969,ProductNode_POSIT4760Output_5892,ProductNode_POSIT4825Output_5970);

SumNode_POSIT1145: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT4825Output_5970,ProductNode_POSIT4721Output_5842,SumNode_POSIT1145Output_5971);

ProductNode_POSIT4826: entity work.PositMult_23_6_comb_uid2(arch)
port map(v13,SumNode_POSIT1145Output_5971,ProductNode_POSIT4826Output_5972);

ProductNode_POSIT4865: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1156Output_6021,ProductNode_POSIT4409Output_5456,ProductNode_POSIT4865Output_6022);

ProductNode_POSIT4897: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT363Output_1901,ProductNode_POSIT4679Output_5790,ProductNode_POSIT4897Output_6060);

ProductNode_POSIT4929: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT369Output_1939,ProductNode_POSIT4711Output_5828,ProductNode_POSIT4929Output_6098);

SumNode_POSIT1169: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT4929Output_6098,ProductNode_POSIT4897Output_6060,SumNode_POSIT1169Output_6099);

ProductNode_POSIT4930: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1169Output_6099,ProductNode_POSIT4865Output_6022,ProductNode_POSIT4930Output_6100);

ProductNode_POSIT4969: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1180Output_6149,ProductNode_POSIT4513Output_5584,ProductNode_POSIT4969Output_6150);

ProductNode_POSIT5001: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT387Output_2029,ProductNode_POSIT4783Output_5918,ProductNode_POSIT5001Output_6188);

ProductNode_POSIT5033: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT393Output_2067,ProductNode_POSIT4815Output_5956,ProductNode_POSIT5033Output_6226);

SumNode_POSIT1193: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT5033Output_6226,ProductNode_POSIT5001Output_6188,SumNode_POSIT1193Output_6227);

ProductNode_POSIT5034: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1193Output_6227,ProductNode_POSIT4969Output_6150,ProductNode_POSIT5034Output_6228);

SumNode_POSIT1194: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT5034Output_6228,ProductNode_POSIT4930Output_6100,SumNode_POSIT1194Output_6229);

ProductNode_POSIT5035: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb13,SumNode_POSIT1194Output_6229,ProductNode_POSIT5035Output_6230);

SumNode_POSIT1195: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT5035Output_6230,ProductNode_POSIT4826Output_5972,SumNode_POSIT1195Output_6231);

ProductNode_POSIT5036: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb3,SumNode_POSIT1195Output_6231,ProductNode_POSIT5036Output_6232);

SumNode_POSIT1196: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT5036Output_6232,ProductNode_POSIT4617Output_5714,SumNode_POSIT1196Output_6233);

ProductNode_POSIT5037: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb4,SumNode_POSIT1196Output_6233,ProductNode_POSIT5037Output_6234);

SumNode_POSIT1197: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT5037Output_6234,ProductNode_POSIT4198Output_5196,SumNode_POSIT1197Output_6235);

ProductNode_POSIT5038: entity work.PositMult_23_6_comb_uid2(arch)
port map(v12,SumNode_POSIT1197Output_6235,ProductNode_POSIT5038Output_6236);

ProductNode_POSIT5040: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT5040weight,ProductNode_POSIT1680Output_2079,ProductNode_POSIT5040Output_6238);

ProductNode_POSIT5042: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT5042weight,v7,ProductNode_POSIT5042Output_6240);

ProductNode_POSIT5043: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT5043weight,vb7,ProductNode_POSIT5043Output_6241);

SumNode_POSIT1198: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT5043Output_6241,ProductNode_POSIT5042Output_6240,SumNode_POSIT1198Output_6242);

ProductNode_POSIT5044: entity work.PositMult_23_6_comb_uid2(arch)
port map(v1,SumNode_POSIT1198Output_6242,ProductNode_POSIT5044Output_6243);

ProductNode_POSIT5049: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1199Output_6248,ProductNode_POSIT5044Output_6243,ProductNode_POSIT5049Output_6249);

ProductNode_POSIT5050: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT5050weight,v7,ProductNode_POSIT5050Output_6250);

ProductNode_POSIT5051: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT5051weight,vb7,ProductNode_POSIT5051Output_6251);

SumNode_POSIT1200: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT5051Output_6251,ProductNode_POSIT5050Output_6250,SumNode_POSIT1200Output_6252);

ProductNode_POSIT5052: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb1,SumNode_POSIT1200Output_6252,ProductNode_POSIT5052Output_6253);

ProductNode_POSIT5057: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1201Output_6258,ProductNode_POSIT5052Output_6253,ProductNode_POSIT5057Output_6259);

SumNode_POSIT1202: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT5057Output_6259,ProductNode_POSIT5049Output_6249,SumNode_POSIT1202Output_6260);

ProductNode_POSIT5058: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1202Output_6260,ProductNode_POSIT1682Output_2081,ProductNode_POSIT5058Output_6261);

ProductNode_POSIT5067: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT405Output_2113,ProductNode_POSIT5044Output_6243,ProductNode_POSIT5067Output_6272);

ProductNode_POSIT5075: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT407Output_2123,ProductNode_POSIT5052Output_6253,ProductNode_POSIT5075Output_6282);

SumNode_POSIT1207: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT5075Output_6282,ProductNode_POSIT5067Output_6272,SumNode_POSIT1207Output_6283);

ProductNode_POSIT5076: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1207Output_6283,ProductNode_POSIT1700Output_2104,ProductNode_POSIT5076Output_6284);

SumNode_POSIT1208: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT5076Output_6284,ProductNode_POSIT5058Output_6261,SumNode_POSIT1208Output_6285);

ProductNode_POSIT5077: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1208Output_6285,ProductNode_POSIT5040Output_6238,ProductNode_POSIT5077Output_6286);

ProductNode_POSIT5109: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT415Output_2165,ProductNode_POSIT3421Output_4234,ProductNode_POSIT5109Output_6324);

ProductNode_POSIT5141: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT421Output_2203,ProductNode_POSIT3453Output_4272,ProductNode_POSIT5141Output_6362);

SumNode_POSIT1221: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT5141Output_6362,ProductNode_POSIT5109Output_6324,SumNode_POSIT1221Output_6363);

ProductNode_POSIT5142: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1221Output_6363,ProductNode_POSIT5077Output_6286,ProductNode_POSIT5142Output_6364);

ProductNode_POSIT5144: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT5144weight,ProductNode_POSIT1784Output_2207,ProductNode_POSIT5144Output_6366);

ProductNode_POSIT5153: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT424Output_2218,ProductNode_POSIT5044Output_6243,ProductNode_POSIT5153Output_6377);

ProductNode_POSIT5161: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT426Output_2228,ProductNode_POSIT5052Output_6253,ProductNode_POSIT5161Output_6387);

SumNode_POSIT1226: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT5161Output_6387,ProductNode_POSIT5153Output_6377,SumNode_POSIT1226Output_6388);

ProductNode_POSIT5162: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1226Output_6388,ProductNode_POSIT1682Output_2081,ProductNode_POSIT5162Output_6389);

ProductNode_POSIT5171: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT429Output_2241,ProductNode_POSIT5044Output_6243,ProductNode_POSIT5171Output_6400);

ProductNode_POSIT5179: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT431Output_2251,ProductNode_POSIT5052Output_6253,ProductNode_POSIT5179Output_6410);

SumNode_POSIT1231: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT5179Output_6410,ProductNode_POSIT5171Output_6400,SumNode_POSIT1231Output_6411);

ProductNode_POSIT5180: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1231Output_6411,ProductNode_POSIT1700Output_2104,ProductNode_POSIT5180Output_6412);

SumNode_POSIT1232: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT5180Output_6412,ProductNode_POSIT5162Output_6389,SumNode_POSIT1232Output_6413);

ProductNode_POSIT5181: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1232Output_6413,ProductNode_POSIT5144Output_6366,ProductNode_POSIT5181Output_6414);

ProductNode_POSIT5213: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT439Output_2293,ProductNode_POSIT3525Output_4362,ProductNode_POSIT5213Output_6452);

ProductNode_POSIT5245: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT445Output_2331,ProductNode_POSIT3557Output_4400,ProductNode_POSIT5245Output_6490);

SumNode_POSIT1245: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT5245Output_6490,ProductNode_POSIT5213Output_6452,SumNode_POSIT1245Output_6491);

ProductNode_POSIT5246: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1245Output_6491,ProductNode_POSIT5181Output_6414,ProductNode_POSIT5246Output_6492);

SumNode_POSIT1246: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT5246Output_6492,ProductNode_POSIT5142Output_6364,SumNode_POSIT1246Output_6493);

ProductNode_POSIT5247: entity work.PositMult_23_6_comb_uid2(arch)
port map(v13,SumNode_POSIT1246Output_6493,ProductNode_POSIT5247Output_6494);

ProductNode_POSIT5249: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT5249weight,ProductNode_POSIT1680Output_2079,ProductNode_POSIT5249Output_6496);

ProductNode_POSIT5286: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1257Output_6543,ProductNode_POSIT5249Output_6496,ProductNode_POSIT5286Output_6544);

ProductNode_POSIT5318: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT464Output_2423,ProductNode_POSIT3421Output_4234,ProductNode_POSIT5318Output_6582);

ProductNode_POSIT5350: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT470Output_2461,ProductNode_POSIT3453Output_4272,ProductNode_POSIT5350Output_6620);

SumNode_POSIT1270: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT5350Output_6620,ProductNode_POSIT5318Output_6582,SumNode_POSIT1270Output_6621);

ProductNode_POSIT5351: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1270Output_6621,ProductNode_POSIT5286Output_6544,ProductNode_POSIT5351Output_6622);

ProductNode_POSIT5353: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT5353weight,ProductNode_POSIT1784Output_2207,ProductNode_POSIT5353Output_6624);

ProductNode_POSIT5390: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1281Output_6671,ProductNode_POSIT5353Output_6624,ProductNode_POSIT5390Output_6672);

ProductNode_POSIT5422: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT488Output_2551,ProductNode_POSIT3525Output_4362,ProductNode_POSIT5422Output_6710);

ProductNode_POSIT5454: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT494Output_2589,ProductNode_POSIT3557Output_4400,ProductNode_POSIT5454Output_6748);

SumNode_POSIT1294: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT5454Output_6748,ProductNode_POSIT5422Output_6710,SumNode_POSIT1294Output_6749);

ProductNode_POSIT5455: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1294Output_6749,ProductNode_POSIT5390Output_6672,ProductNode_POSIT5455Output_6750);

SumNode_POSIT1295: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT5455Output_6750,ProductNode_POSIT5351Output_6622,SumNode_POSIT1295Output_6751);

ProductNode_POSIT5456: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb13,SumNode_POSIT1295Output_6751,ProductNode_POSIT5456Output_6752);

SumNode_POSIT1296: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT5456Output_6752,ProductNode_POSIT5247Output_6494,SumNode_POSIT1296Output_6753);

ProductNode_POSIT5457: entity work.PositMult_23_6_comb_uid2(arch)
port map(v3,SumNode_POSIT1296Output_6753,ProductNode_POSIT5457Output_6754);

ProductNode_POSIT5477: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1301Output_6778,ProductNode_POSIT2101Output_2599,ProductNode_POSIT5477Output_6779);

ProductNode_POSIT5495: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1306Output_6801,ProductNode_POSIT2119Output_2622,ProductNode_POSIT5495Output_6802);

SumNode_POSIT1307: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT5495Output_6802,ProductNode_POSIT5477Output_6779,SumNode_POSIT1307Output_6803);

ProductNode_POSIT5496: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1307Output_6803,ProductNode_POSIT5040Output_6238,ProductNode_POSIT5496Output_6804);

ProductNode_POSIT5528: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT514Output_2683,ProductNode_POSIT3840Output_4752,ProductNode_POSIT5528Output_6842);

ProductNode_POSIT5560: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT520Output_2721,ProductNode_POSIT3872Output_4790,ProductNode_POSIT5560Output_6880);

SumNode_POSIT1320: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT5560Output_6880,ProductNode_POSIT5528Output_6842,SumNode_POSIT1320Output_6881);

ProductNode_POSIT5561: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1320Output_6881,ProductNode_POSIT5496Output_6804,ProductNode_POSIT5561Output_6882);

ProductNode_POSIT5581: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1325Output_6906,ProductNode_POSIT2101Output_2599,ProductNode_POSIT5581Output_6907);

ProductNode_POSIT5599: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1330Output_6929,ProductNode_POSIT2119Output_2622,ProductNode_POSIT5599Output_6930);

SumNode_POSIT1331: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT5599Output_6930,ProductNode_POSIT5581Output_6907,SumNode_POSIT1331Output_6931);

ProductNode_POSIT5600: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1331Output_6931,ProductNode_POSIT5144Output_6366,ProductNode_POSIT5600Output_6932);

ProductNode_POSIT5632: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT538Output_2811,ProductNode_POSIT3944Output_4880,ProductNode_POSIT5632Output_6970);

ProductNode_POSIT5664: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT544Output_2849,ProductNode_POSIT3976Output_4918,ProductNode_POSIT5664Output_7008);

SumNode_POSIT1344: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT5664Output_7008,ProductNode_POSIT5632Output_6970,SumNode_POSIT1344Output_7009);

ProductNode_POSIT5665: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1344Output_7009,ProductNode_POSIT5600Output_6932,ProductNode_POSIT5665Output_7010);

SumNode_POSIT1345: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT5665Output_7010,ProductNode_POSIT5561Output_6882,SumNode_POSIT1345Output_7011);

ProductNode_POSIT5666: entity work.PositMult_23_6_comb_uid2(arch)
port map(v13,SumNode_POSIT1345Output_7011,ProductNode_POSIT5666Output_7012);

ProductNode_POSIT5705: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1356Output_7061,ProductNode_POSIT5249Output_6496,ProductNode_POSIT5705Output_7062);

ProductNode_POSIT5737: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT563Output_2941,ProductNode_POSIT3840Output_4752,ProductNode_POSIT5737Output_7100);

ProductNode_POSIT5769: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT569Output_2979,ProductNode_POSIT3872Output_4790,ProductNode_POSIT5769Output_7138);

SumNode_POSIT1369: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT5769Output_7138,ProductNode_POSIT5737Output_7100,SumNode_POSIT1369Output_7139);

ProductNode_POSIT5770: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1369Output_7139,ProductNode_POSIT5705Output_7062,ProductNode_POSIT5770Output_7140);

ProductNode_POSIT5809: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1380Output_7189,ProductNode_POSIT5353Output_6624,ProductNode_POSIT5809Output_7190);

ProductNode_POSIT5841: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT587Output_3069,ProductNode_POSIT3944Output_4880,ProductNode_POSIT5841Output_7228);

ProductNode_POSIT5873: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT593Output_3107,ProductNode_POSIT3976Output_4918,ProductNode_POSIT5873Output_7266);

SumNode_POSIT1393: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT5873Output_7266,ProductNode_POSIT5841Output_7228,SumNode_POSIT1393Output_7267);

ProductNode_POSIT5874: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1393Output_7267,ProductNode_POSIT5809Output_7190,ProductNode_POSIT5874Output_7268);

SumNode_POSIT1394: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT5874Output_7268,ProductNode_POSIT5770Output_7140,SumNode_POSIT1394Output_7269);

ProductNode_POSIT5875: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb13,SumNode_POSIT1394Output_7269,ProductNode_POSIT5875Output_7270);

SumNode_POSIT1395: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT5875Output_7270,ProductNode_POSIT5666Output_7012,SumNode_POSIT1395Output_7271);

ProductNode_POSIT5876: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb3,SumNode_POSIT1395Output_7271,ProductNode_POSIT5876Output_7272);

SumNode_POSIT1396: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT5876Output_7272,ProductNode_POSIT5457Output_6754,SumNode_POSIT1396Output_7273);

ProductNode_POSIT5877: entity work.PositMult_23_6_comb_uid2(arch)
port map(v4,SumNode_POSIT1396Output_7273,ProductNode_POSIT5877Output_7274);

ProductNode_POSIT5879: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT5879weight,ProductNode_POSIT2519Output_3117,ProductNode_POSIT5879Output_7276);

ProductNode_POSIT5881: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT5881weight,v7,ProductNode_POSIT5881Output_7278);

ProductNode_POSIT5882: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT5882weight,vb7,ProductNode_POSIT5882Output_7279);

SumNode_POSIT1397: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT5882Output_7279,ProductNode_POSIT5881Output_7278,SumNode_POSIT1397Output_7280);

ProductNode_POSIT5883: entity work.PositMult_23_6_comb_uid2(arch)
port map(v1,SumNode_POSIT1397Output_7280,ProductNode_POSIT5883Output_7281);

ProductNode_POSIT5888: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1398Output_7286,ProductNode_POSIT5883Output_7281,ProductNode_POSIT5888Output_7287);

ProductNode_POSIT5889: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT5889weight,v7,ProductNode_POSIT5889Output_7288);

ProductNode_POSIT5890: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT5890weight,vb7,ProductNode_POSIT5890Output_7289);

SumNode_POSIT1399: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT5890Output_7289,ProductNode_POSIT5889Output_7288,SumNode_POSIT1399Output_7290);

ProductNode_POSIT5891: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb1,SumNode_POSIT1399Output_7290,ProductNode_POSIT5891Output_7291);

ProductNode_POSIT5896: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1400Output_7296,ProductNode_POSIT5891Output_7291,ProductNode_POSIT5896Output_7297);

SumNode_POSIT1401: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT5896Output_7297,ProductNode_POSIT5888Output_7287,SumNode_POSIT1401Output_7298);

ProductNode_POSIT5897: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1401Output_7298,ProductNode_POSIT2521Output_3119,ProductNode_POSIT5897Output_7299);

ProductNode_POSIT5906: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT405Output_2113,ProductNode_POSIT5883Output_7281,ProductNode_POSIT5906Output_7310);

ProductNode_POSIT5914: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT407Output_2123,ProductNode_POSIT5891Output_7291,ProductNode_POSIT5914Output_7320);

SumNode_POSIT1406: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT5914Output_7320,ProductNode_POSIT5906Output_7310,SumNode_POSIT1406Output_7321);

ProductNode_POSIT5915: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1406Output_7321,ProductNode_POSIT2539Output_3142,ProductNode_POSIT5915Output_7322);

SumNode_POSIT1407: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT5915Output_7322,ProductNode_POSIT5897Output_7299,SumNode_POSIT1407Output_7323);

ProductNode_POSIT5916: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1407Output_7323,ProductNode_POSIT5879Output_7276,ProductNode_POSIT5916Output_7324);

ProductNode_POSIT5948: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT614Output_3203,ProductNode_POSIT4260Output_5272,ProductNode_POSIT5948Output_7362);

ProductNode_POSIT5980: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT620Output_3241,ProductNode_POSIT4292Output_5310,ProductNode_POSIT5980Output_7400);

SumNode_POSIT1420: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT5980Output_7400,ProductNode_POSIT5948Output_7362,SumNode_POSIT1420Output_7401);

ProductNode_POSIT5981: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1420Output_7401,ProductNode_POSIT5916Output_7324,ProductNode_POSIT5981Output_7402);

ProductNode_POSIT5983: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT5983weight,ProductNode_POSIT2623Output_3245,ProductNode_POSIT5983Output_7404);

ProductNode_POSIT5992: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT424Output_2218,ProductNode_POSIT5883Output_7281,ProductNode_POSIT5992Output_7415);

ProductNode_POSIT6000: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT426Output_2228,ProductNode_POSIT5891Output_7291,ProductNode_POSIT6000Output_7425);

SumNode_POSIT1425: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT6000Output_7425,ProductNode_POSIT5992Output_7415,SumNode_POSIT1425Output_7426);

ProductNode_POSIT6001: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1425Output_7426,ProductNode_POSIT2521Output_3119,ProductNode_POSIT6001Output_7427);

ProductNode_POSIT6010: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT429Output_2241,ProductNode_POSIT5883Output_7281,ProductNode_POSIT6010Output_7438);

ProductNode_POSIT6018: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT431Output_2251,ProductNode_POSIT5891Output_7291,ProductNode_POSIT6018Output_7448);

SumNode_POSIT1430: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT6018Output_7448,ProductNode_POSIT6010Output_7438,SumNode_POSIT1430Output_7449);

ProductNode_POSIT6019: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1430Output_7449,ProductNode_POSIT2539Output_3142,ProductNode_POSIT6019Output_7450);

SumNode_POSIT1431: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT6019Output_7450,ProductNode_POSIT6001Output_7427,SumNode_POSIT1431Output_7451);

ProductNode_POSIT6020: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1431Output_7451,ProductNode_POSIT5983Output_7404,ProductNode_POSIT6020Output_7452);

ProductNode_POSIT6052: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT638Output_3331,ProductNode_POSIT4364Output_5400,ProductNode_POSIT6052Output_7490);

ProductNode_POSIT6084: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT644Output_3369,ProductNode_POSIT4396Output_5438,ProductNode_POSIT6084Output_7528);

SumNode_POSIT1444: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT6084Output_7528,ProductNode_POSIT6052Output_7490,SumNode_POSIT1444Output_7529);

ProductNode_POSIT6085: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1444Output_7529,ProductNode_POSIT6020Output_7452,ProductNode_POSIT6085Output_7530);

SumNode_POSIT1445: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT6085Output_7530,ProductNode_POSIT5981Output_7402,SumNode_POSIT1445Output_7531);

ProductNode_POSIT6086: entity work.PositMult_23_6_comb_uid2(arch)
port map(v13,SumNode_POSIT1445Output_7531,ProductNode_POSIT6086Output_7532);

ProductNode_POSIT6088: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT6088weight,ProductNode_POSIT2519Output_3117,ProductNode_POSIT6088Output_7534);

ProductNode_POSIT6125: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1456Output_7581,ProductNode_POSIT6088Output_7534,ProductNode_POSIT6125Output_7582);

ProductNode_POSIT6157: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT663Output_3461,ProductNode_POSIT4260Output_5272,ProductNode_POSIT6157Output_7620);

ProductNode_POSIT6189: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT669Output_3499,ProductNode_POSIT4292Output_5310,ProductNode_POSIT6189Output_7658);

SumNode_POSIT1469: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT6189Output_7658,ProductNode_POSIT6157Output_7620,SumNode_POSIT1469Output_7659);

ProductNode_POSIT6190: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1469Output_7659,ProductNode_POSIT6125Output_7582,ProductNode_POSIT6190Output_7660);

ProductNode_POSIT6192: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT6192weight,ProductNode_POSIT2623Output_3245,ProductNode_POSIT6192Output_7662);

ProductNode_POSIT6229: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1480Output_7709,ProductNode_POSIT6192Output_7662,ProductNode_POSIT6229Output_7710);

ProductNode_POSIT6261: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT687Output_3589,ProductNode_POSIT4364Output_5400,ProductNode_POSIT6261Output_7748);

ProductNode_POSIT6293: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT693Output_3627,ProductNode_POSIT4396Output_5438,ProductNode_POSIT6293Output_7786);

SumNode_POSIT1493: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT6293Output_7786,ProductNode_POSIT6261Output_7748,SumNode_POSIT1493Output_7787);

ProductNode_POSIT6294: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1493Output_7787,ProductNode_POSIT6229Output_7710,ProductNode_POSIT6294Output_7788);

SumNode_POSIT1494: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT6294Output_7788,ProductNode_POSIT6190Output_7660,SumNode_POSIT1494Output_7789);

ProductNode_POSIT6295: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb13,SumNode_POSIT1494Output_7789,ProductNode_POSIT6295Output_7790);

SumNode_POSIT1495: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT6295Output_7790,ProductNode_POSIT6086Output_7532,SumNode_POSIT1495Output_7791);

ProductNode_POSIT6296: entity work.PositMult_23_6_comb_uid2(arch)
port map(v3,SumNode_POSIT1495Output_7791,ProductNode_POSIT6296Output_7792);

ProductNode_POSIT6316: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1500Output_7816,ProductNode_POSIT2940Output_3637,ProductNode_POSIT6316Output_7817);

ProductNode_POSIT6334: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1505Output_7839,ProductNode_POSIT2958Output_3660,ProductNode_POSIT6334Output_7840);

SumNode_POSIT1506: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT6334Output_7840,ProductNode_POSIT6316Output_7817,SumNode_POSIT1506Output_7841);

ProductNode_POSIT6335: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1506Output_7841,ProductNode_POSIT5879Output_7276,ProductNode_POSIT6335Output_7842);

ProductNode_POSIT6367: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT713Output_3721,ProductNode_POSIT4679Output_5790,ProductNode_POSIT6367Output_7880);

ProductNode_POSIT6399: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT719Output_3759,ProductNode_POSIT4711Output_5828,ProductNode_POSIT6399Output_7918);

SumNode_POSIT1519: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT6399Output_7918,ProductNode_POSIT6367Output_7880,SumNode_POSIT1519Output_7919);

ProductNode_POSIT6400: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1519Output_7919,ProductNode_POSIT6335Output_7842,ProductNode_POSIT6400Output_7920);

ProductNode_POSIT6420: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1524Output_7944,ProductNode_POSIT2940Output_3637,ProductNode_POSIT6420Output_7945);

ProductNode_POSIT6438: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1529Output_7967,ProductNode_POSIT2958Output_3660,ProductNode_POSIT6438Output_7968);

SumNode_POSIT1530: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT6438Output_7968,ProductNode_POSIT6420Output_7945,SumNode_POSIT1530Output_7969);

ProductNode_POSIT6439: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1530Output_7969,ProductNode_POSIT5983Output_7404,ProductNode_POSIT6439Output_7970);

ProductNode_POSIT6471: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT737Output_3849,ProductNode_POSIT4783Output_5918,ProductNode_POSIT6471Output_8008);

ProductNode_POSIT6503: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT743Output_3887,ProductNode_POSIT4815Output_5956,ProductNode_POSIT6503Output_8046);

SumNode_POSIT1543: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT6503Output_8046,ProductNode_POSIT6471Output_8008,SumNode_POSIT1543Output_8047);

ProductNode_POSIT6504: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1543Output_8047,ProductNode_POSIT6439Output_7970,ProductNode_POSIT6504Output_8048);

SumNode_POSIT1544: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT6504Output_8048,ProductNode_POSIT6400Output_7920,SumNode_POSIT1544Output_8049);

ProductNode_POSIT6505: entity work.PositMult_23_6_comb_uid2(arch)
port map(v13,SumNode_POSIT1544Output_8049,ProductNode_POSIT6505Output_8050);

ProductNode_POSIT6544: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1555Output_8099,ProductNode_POSIT6088Output_7534,ProductNode_POSIT6544Output_8100);

ProductNode_POSIT6576: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT762Output_3979,ProductNode_POSIT4679Output_5790,ProductNode_POSIT6576Output_8138);

ProductNode_POSIT6608: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT768Output_4017,ProductNode_POSIT4711Output_5828,ProductNode_POSIT6608Output_8176);

SumNode_POSIT1568: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT6608Output_8176,ProductNode_POSIT6576Output_8138,SumNode_POSIT1568Output_8177);

ProductNode_POSIT6609: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1568Output_8177,ProductNode_POSIT6544Output_8100,ProductNode_POSIT6609Output_8178);

ProductNode_POSIT6648: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1579Output_8227,ProductNode_POSIT6192Output_7662,ProductNode_POSIT6648Output_8228);

ProductNode_POSIT6680: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT786Output_4107,ProductNode_POSIT4783Output_5918,ProductNode_POSIT6680Output_8266);

ProductNode_POSIT6712: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT792Output_4145,ProductNode_POSIT4815Output_5956,ProductNode_POSIT6712Output_8304);

SumNode_POSIT1592: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT6712Output_8304,ProductNode_POSIT6680Output_8266,SumNode_POSIT1592Output_8305);

ProductNode_POSIT6713: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1592Output_8305,ProductNode_POSIT6648Output_8228,ProductNode_POSIT6713Output_8306);

SumNode_POSIT1593: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT6713Output_8306,ProductNode_POSIT6609Output_8178,SumNode_POSIT1593Output_8307);

ProductNode_POSIT6714: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb13,SumNode_POSIT1593Output_8307,ProductNode_POSIT6714Output_8308);

SumNode_POSIT1594: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT6714Output_8308,ProductNode_POSIT6505Output_8050,SumNode_POSIT1594Output_8309);

ProductNode_POSIT6715: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb3,SumNode_POSIT1594Output_8309,ProductNode_POSIT6715Output_8310);

SumNode_POSIT1595: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT6715Output_8310,ProductNode_POSIT6296Output_7792,SumNode_POSIT1595Output_8311);

ProductNode_POSIT6716: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb4,SumNode_POSIT1595Output_8311,ProductNode_POSIT6716Output_8312);

SumNode_POSIT1596: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT6716Output_8312,ProductNode_POSIT5877Output_7274,SumNode_POSIT1596Output_8313);

ProductNode_POSIT6717: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb12,SumNode_POSIT1596Output_8313,ProductNode_POSIT6717Output_8314);

SumNode_POSIT1597: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT6717Output_8314,ProductNode_POSIT5038Output_6236,SumNode_POSIT1597Output_8315);

ProductNode_POSIT6718: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb6,SumNode_POSIT1597Output_8315,ProductNode_POSIT6718Output_8316);

SumNode_POSIT1598: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT6718Output_8316,ProductNode_POSIT3359Output_4158,SumNode_POSIT1598Output_8317);

ProductNode_POSIT6719: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1598Output_8317,ProductNode_POSIT0Output_0,ProductNode_POSIT6719Output_8318);

ProductNode_POSIT6720: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT6720weight,vb9,ProductNode_POSIT6720Output_8319);

ProductNode_POSIT6722: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT6722weight,ProductNode_POSIT1Output_1,ProductNode_POSIT6722Output_8321);

ProductNode_POSIT6728: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT6728weight,ProductNode_POSIT7Output_8,ProductNode_POSIT6728Output_8328);

ProductNode_POSIT6730: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT6730weight,ProductNode_POSIT9Output_10,ProductNode_POSIT6730Output_8330);

SumNode_POSIT1600: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT6730Output_8330,ProductNode_POSIT6728Output_8328,SumNode_POSIT1600Output_8331);

ProductNode_POSIT6731: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1600Output_8331,ProductNode_POSIT6Output_7,ProductNode_POSIT6731Output_8332);

ProductNode_POSIT6736: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT6736weight,ProductNode_POSIT15Output_18,ProductNode_POSIT6736Output_8338);

ProductNode_POSIT6738: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT6738weight,ProductNode_POSIT17Output_20,ProductNode_POSIT6738Output_8340);

SumNode_POSIT1602: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT6738Output_8340,ProductNode_POSIT6736Output_8338,SumNode_POSIT1602Output_8341);

ProductNode_POSIT6739: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1602Output_8341,ProductNode_POSIT14Output_17,ProductNode_POSIT6739Output_8342);

SumNode_POSIT1603: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT6739Output_8342,ProductNode_POSIT6731Output_8332,SumNode_POSIT1603Output_8343);

ProductNode_POSIT6740: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1603Output_8343,ProductNode_POSIT3Output_3,ProductNode_POSIT6740Output_8344);

ProductNode_POSIT6746: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT6746weight,ProductNode_POSIT25Output_31,ProductNode_POSIT6746Output_8351);

ProductNode_POSIT6748: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT6748weight,ProductNode_POSIT27Output_33,ProductNode_POSIT6748Output_8353);

SumNode_POSIT1605: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT6748Output_8353,ProductNode_POSIT6746Output_8351,SumNode_POSIT1605Output_8354);

ProductNode_POSIT6749: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1605Output_8354,ProductNode_POSIT6Output_7,ProductNode_POSIT6749Output_8355);

ProductNode_POSIT6754: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT6754weight,ProductNode_POSIT33Output_41,ProductNode_POSIT6754Output_8361);

ProductNode_POSIT6756: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT6756weight,ProductNode_POSIT35Output_43,ProductNode_POSIT6756Output_8363);

SumNode_POSIT1607: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT6756Output_8363,ProductNode_POSIT6754Output_8361,SumNode_POSIT1607Output_8364);

ProductNode_POSIT6757: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1607Output_8364,ProductNode_POSIT14Output_17,ProductNode_POSIT6757Output_8365);

SumNode_POSIT1608: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT6757Output_8365,ProductNode_POSIT6749Output_8355,SumNode_POSIT1608Output_8366);

ProductNode_POSIT6758: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1608Output_8366,ProductNode_POSIT21Output_26,ProductNode_POSIT6758Output_8367);

SumNode_POSIT1609: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT6758Output_8367,ProductNode_POSIT6740Output_8344,SumNode_POSIT1609Output_8368);

ProductNode_POSIT6759: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1609Output_8368,ProductNode_POSIT6722Output_8321,ProductNode_POSIT6759Output_8369);

ProductNode_POSIT6760: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT6760weight,v10,ProductNode_POSIT6760Output_8370);

ProductNode_POSIT6781: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1612Output_8393,ProductNode_POSIT6760Output_8370,ProductNode_POSIT6781Output_8394);

ProductNode_POSIT6782: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT6782weight,ProductNode_POSIT6781Output_8394,ProductNode_POSIT6782Output_8395);

ProductNode_POSIT6786: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT6786weight,ProductNode_POSIT65Output_80,ProductNode_POSIT6786Output_8400);

ProductNode_POSIT6790: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT6790weight,ProductNode_POSIT69Output_85,ProductNode_POSIT6790Output_8405);

SumNode_POSIT1615: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT6790Output_8405,ProductNode_POSIT6786Output_8400,SumNode_POSIT1615Output_8406);

ProductNode_POSIT6791: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1615Output_8406,ProductNode_POSIT6782Output_8395,ProductNode_POSIT6791Output_8407);

ProductNode_POSIT6792: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT6792weight,vb10,ProductNode_POSIT6792Output_8408);

ProductNode_POSIT6813: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1618Output_8431,ProductNode_POSIT6792Output_8408,ProductNode_POSIT6813Output_8432);

ProductNode_POSIT6814: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT6814weight,ProductNode_POSIT6813Output_8432,ProductNode_POSIT6814Output_8433);

ProductNode_POSIT6818: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT6818weight,ProductNode_POSIT65Output_80,ProductNode_POSIT6818Output_8438);

ProductNode_POSIT6822: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT6822weight,ProductNode_POSIT69Output_85,ProductNode_POSIT6822Output_8443);

SumNode_POSIT1621: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT6822Output_8443,ProductNode_POSIT6818Output_8438,SumNode_POSIT1621Output_8444);

ProductNode_POSIT6823: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1621Output_8444,ProductNode_POSIT6814Output_8433,ProductNode_POSIT6823Output_8445);

SumNode_POSIT1622: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT6823Output_8445,ProductNode_POSIT6791Output_8407,SumNode_POSIT1622Output_8446);

ProductNode_POSIT6824: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1622Output_8446,ProductNode_POSIT6759Output_8369,ProductNode_POSIT6824Output_8447);

ProductNode_POSIT6826: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT6826weight,ProductNode_POSIT105Output_129,ProductNode_POSIT6826Output_8449);

ProductNode_POSIT6832: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT6832weight,ProductNode_POSIT7Output_8,ProductNode_POSIT6832Output_8456);

ProductNode_POSIT6834: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT6834weight,ProductNode_POSIT9Output_10,ProductNode_POSIT6834Output_8458);

SumNode_POSIT1624: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT6834Output_8458,ProductNode_POSIT6832Output_8456,SumNode_POSIT1624Output_8459);

ProductNode_POSIT6835: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1624Output_8459,ProductNode_POSIT6Output_7,ProductNode_POSIT6835Output_8460);

ProductNode_POSIT6840: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT6840weight,ProductNode_POSIT15Output_18,ProductNode_POSIT6840Output_8466);

ProductNode_POSIT6842: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT6842weight,ProductNode_POSIT17Output_20,ProductNode_POSIT6842Output_8468);

SumNode_POSIT1626: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT6842Output_8468,ProductNode_POSIT6840Output_8466,SumNode_POSIT1626Output_8469);

ProductNode_POSIT6843: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1626Output_8469,ProductNode_POSIT14Output_17,ProductNode_POSIT6843Output_8470);

SumNode_POSIT1627: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT6843Output_8470,ProductNode_POSIT6835Output_8460,SumNode_POSIT1627Output_8471);

ProductNode_POSIT6844: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1627Output_8471,ProductNode_POSIT3Output_3,ProductNode_POSIT6844Output_8472);

ProductNode_POSIT6850: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT6850weight,ProductNode_POSIT25Output_31,ProductNode_POSIT6850Output_8479);

ProductNode_POSIT6852: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT6852weight,ProductNode_POSIT27Output_33,ProductNode_POSIT6852Output_8481);

SumNode_POSIT1629: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT6852Output_8481,ProductNode_POSIT6850Output_8479,SumNode_POSIT1629Output_8482);

ProductNode_POSIT6853: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1629Output_8482,ProductNode_POSIT6Output_7,ProductNode_POSIT6853Output_8483);

ProductNode_POSIT6858: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT6858weight,ProductNode_POSIT33Output_41,ProductNode_POSIT6858Output_8489);

ProductNode_POSIT6860: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT6860weight,ProductNode_POSIT35Output_43,ProductNode_POSIT6860Output_8491);

SumNode_POSIT1631: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT6860Output_8491,ProductNode_POSIT6858Output_8489,SumNode_POSIT1631Output_8492);

ProductNode_POSIT6861: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1631Output_8492,ProductNode_POSIT14Output_17,ProductNode_POSIT6861Output_8493);

SumNode_POSIT1632: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT6861Output_8493,ProductNode_POSIT6853Output_8483,SumNode_POSIT1632Output_8494);

ProductNode_POSIT6862: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1632Output_8494,ProductNode_POSIT21Output_26,ProductNode_POSIT6862Output_8495);

SumNode_POSIT1633: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT6862Output_8495,ProductNode_POSIT6844Output_8472,SumNode_POSIT1633Output_8496);

ProductNode_POSIT6863: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1633Output_8496,ProductNode_POSIT6826Output_8449,ProductNode_POSIT6863Output_8497);

ProductNode_POSIT6886: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT6886weight,ProductNode_POSIT6781Output_8394,ProductNode_POSIT6886Output_8523);

ProductNode_POSIT6890: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT6890weight,ProductNode_POSIT65Output_80,ProductNode_POSIT6890Output_8528);

ProductNode_POSIT6894: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT6894weight,ProductNode_POSIT69Output_85,ProductNode_POSIT6894Output_8533);

SumNode_POSIT1639: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT6894Output_8533,ProductNode_POSIT6890Output_8528,SumNode_POSIT1639Output_8534);

ProductNode_POSIT6895: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1639Output_8534,ProductNode_POSIT6886Output_8523,ProductNode_POSIT6895Output_8535);

ProductNode_POSIT6918: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT6918weight,ProductNode_POSIT6813Output_8432,ProductNode_POSIT6918Output_8561);

ProductNode_POSIT6922: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT6922weight,ProductNode_POSIT65Output_80,ProductNode_POSIT6922Output_8566);

ProductNode_POSIT6926: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT6926weight,ProductNode_POSIT69Output_85,ProductNode_POSIT6926Output_8571);

SumNode_POSIT1645: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT6926Output_8571,ProductNode_POSIT6922Output_8566,SumNode_POSIT1645Output_8572);

ProductNode_POSIT6927: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1645Output_8572,ProductNode_POSIT6918Output_8561,ProductNode_POSIT6927Output_8573);

SumNode_POSIT1646: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT6927Output_8573,ProductNode_POSIT6895Output_8535,SumNode_POSIT1646Output_8574);

ProductNode_POSIT6928: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1646Output_8574,ProductNode_POSIT6863Output_8497,ProductNode_POSIT6928Output_8575);

SumNode_POSIT1647: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT6928Output_8575,ProductNode_POSIT6824Output_8447,SumNode_POSIT1647Output_8576);

ProductNode_POSIT6929: entity work.PositMult_23_6_comb_uid2(arch)
port map(v13,SumNode_POSIT1647Output_8576,ProductNode_POSIT6929Output_8577);

ProductNode_POSIT6931: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT6931weight,ProductNode_POSIT1Output_1,ProductNode_POSIT6931Output_8579);

ProductNode_POSIT6968: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1658Output_8626,ProductNode_POSIT6931Output_8579,ProductNode_POSIT6968Output_8627);

ProductNode_POSIT6995: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT6995weight,ProductNode_POSIT274Output_338,ProductNode_POSIT6995Output_8658);

ProductNode_POSIT6999: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT6999weight,ProductNode_POSIT278Output_343,ProductNode_POSIT6999Output_8663);

SumNode_POSIT1664: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT6999Output_8663,ProductNode_POSIT6995Output_8658,SumNode_POSIT1664Output_8664);

ProductNode_POSIT7000: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1664Output_8664,ProductNode_POSIT6782Output_8395,ProductNode_POSIT7000Output_8665);

ProductNode_POSIT7027: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT7027weight,ProductNode_POSIT274Output_338,ProductNode_POSIT7027Output_8696);

ProductNode_POSIT7031: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT7031weight,ProductNode_POSIT278Output_343,ProductNode_POSIT7031Output_8701);

SumNode_POSIT1670: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT7031Output_8701,ProductNode_POSIT7027Output_8696,SumNode_POSIT1670Output_8702);

ProductNode_POSIT7032: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1670Output_8702,ProductNode_POSIT6814Output_8433,ProductNode_POSIT7032Output_8703);

SumNode_POSIT1671: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT7032Output_8703,ProductNode_POSIT7000Output_8665,SumNode_POSIT1671Output_8704);

ProductNode_POSIT7033: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1671Output_8704,ProductNode_POSIT6968Output_8627,ProductNode_POSIT7033Output_8705);

ProductNode_POSIT7035: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT7035weight,ProductNode_POSIT105Output_129,ProductNode_POSIT7035Output_8707);

ProductNode_POSIT7072: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1682Output_8754,ProductNode_POSIT7035Output_8707,ProductNode_POSIT7072Output_8755);

ProductNode_POSIT7099: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT7099weight,ProductNode_POSIT274Output_338,ProductNode_POSIT7099Output_8786);

ProductNode_POSIT7103: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT7103weight,ProductNode_POSIT278Output_343,ProductNode_POSIT7103Output_8791);

SumNode_POSIT1688: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT7103Output_8791,ProductNode_POSIT7099Output_8786,SumNode_POSIT1688Output_8792);

ProductNode_POSIT7104: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1688Output_8792,ProductNode_POSIT6886Output_8523,ProductNode_POSIT7104Output_8793);

ProductNode_POSIT7131: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT7131weight,ProductNode_POSIT274Output_338,ProductNode_POSIT7131Output_8824);

ProductNode_POSIT7135: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT7135weight,ProductNode_POSIT278Output_343,ProductNode_POSIT7135Output_8829);

SumNode_POSIT1694: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT7135Output_8829,ProductNode_POSIT7131Output_8824,SumNode_POSIT1694Output_8830);

ProductNode_POSIT7136: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1694Output_8830,ProductNode_POSIT6918Output_8561,ProductNode_POSIT7136Output_8831);

SumNode_POSIT1695: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT7136Output_8831,ProductNode_POSIT7104Output_8793,SumNode_POSIT1695Output_8832);

ProductNode_POSIT7137: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1695Output_8832,ProductNode_POSIT7072Output_8755,ProductNode_POSIT7137Output_8833);

SumNode_POSIT1696: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT7137Output_8833,ProductNode_POSIT7033Output_8705,SumNode_POSIT1696Output_8834);

ProductNode_POSIT7138: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb13,SumNode_POSIT1696Output_8834,ProductNode_POSIT7138Output_8835);

SumNode_POSIT1697: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT7138Output_8835,ProductNode_POSIT6929Output_8577,SumNode_POSIT1697Output_8836);

ProductNode_POSIT7139: entity work.PositMult_23_6_comb_uid2(arch)
port map(v3,SumNode_POSIT1697Output_8836,ProductNode_POSIT7139Output_8837);

ProductNode_POSIT7159: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1702Output_8861,ProductNode_POSIT422Output_521,ProductNode_POSIT7159Output_8862);

ProductNode_POSIT7177: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1707Output_8884,ProductNode_POSIT440Output_544,ProductNode_POSIT7177Output_8885);

SumNode_POSIT1708: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT7177Output_8885,ProductNode_POSIT7159Output_8862,SumNode_POSIT1708Output_8886);

ProductNode_POSIT7178: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1708Output_8886,ProductNode_POSIT6722Output_8321,ProductNode_POSIT7178Output_8887);

ProductNode_POSIT7200: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT112Output_592,ProductNode_POSIT6760Output_8370,ProductNode_POSIT7200Output_8912);

ProductNode_POSIT7201: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT7201weight,ProductNode_POSIT7200Output_8912,ProductNode_POSIT7201Output_8913);

ProductNode_POSIT7205: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT7205weight,ProductNode_POSIT65Output_80,ProductNode_POSIT7205Output_8918);

ProductNode_POSIT7209: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT7209weight,ProductNode_POSIT69Output_85,ProductNode_POSIT7209Output_8923);

SumNode_POSIT1714: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT7209Output_8923,ProductNode_POSIT7205Output_8918,SumNode_POSIT1714Output_8924);

ProductNode_POSIT7210: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1714Output_8924,ProductNode_POSIT7201Output_8913,ProductNode_POSIT7210Output_8925);

ProductNode_POSIT7232: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT118Output_630,ProductNode_POSIT6792Output_8408,ProductNode_POSIT7232Output_8950);

ProductNode_POSIT7233: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT7233weight,ProductNode_POSIT7232Output_8950,ProductNode_POSIT7233Output_8951);

ProductNode_POSIT7237: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT7237weight,ProductNode_POSIT65Output_80,ProductNode_POSIT7237Output_8956);

ProductNode_POSIT7241: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT7241weight,ProductNode_POSIT69Output_85,ProductNode_POSIT7241Output_8961);

SumNode_POSIT1720: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT7241Output_8961,ProductNode_POSIT7237Output_8956,SumNode_POSIT1720Output_8962);

ProductNode_POSIT7242: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1720Output_8962,ProductNode_POSIT7233Output_8951,ProductNode_POSIT7242Output_8963);

SumNode_POSIT1721: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT7242Output_8963,ProductNode_POSIT7210Output_8925,SumNode_POSIT1721Output_8964);

ProductNode_POSIT7243: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1721Output_8964,ProductNode_POSIT7178Output_8887,ProductNode_POSIT7243Output_8965);

ProductNode_POSIT7263: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1726Output_8989,ProductNode_POSIT422Output_521,ProductNode_POSIT7263Output_8990);

ProductNode_POSIT7281: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1731Output_9012,ProductNode_POSIT440Output_544,ProductNode_POSIT7281Output_9013);

SumNode_POSIT1732: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT7281Output_9013,ProductNode_POSIT7263Output_8990,SumNode_POSIT1732Output_9014);

ProductNode_POSIT7282: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1732Output_9014,ProductNode_POSIT6826Output_8449,ProductNode_POSIT7282Output_9015);

ProductNode_POSIT7305: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT7305weight,ProductNode_POSIT7200Output_8912,ProductNode_POSIT7305Output_9041);

ProductNode_POSIT7309: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT7309weight,ProductNode_POSIT65Output_80,ProductNode_POSIT7309Output_9046);

ProductNode_POSIT7313: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT7313weight,ProductNode_POSIT69Output_85,ProductNode_POSIT7313Output_9051);

SumNode_POSIT1738: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT7313Output_9051,ProductNode_POSIT7309Output_9046,SumNode_POSIT1738Output_9052);

ProductNode_POSIT7314: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1738Output_9052,ProductNode_POSIT7305Output_9041,ProductNode_POSIT7314Output_9053);

ProductNode_POSIT7337: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT7337weight,ProductNode_POSIT7232Output_8950,ProductNode_POSIT7337Output_9079);

ProductNode_POSIT7341: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT7341weight,ProductNode_POSIT65Output_80,ProductNode_POSIT7341Output_9084);

ProductNode_POSIT7345: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT7345weight,ProductNode_POSIT69Output_85,ProductNode_POSIT7345Output_9089);

SumNode_POSIT1744: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT7345Output_9089,ProductNode_POSIT7341Output_9084,SumNode_POSIT1744Output_9090);

ProductNode_POSIT7346: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1744Output_9090,ProductNode_POSIT7337Output_9079,ProductNode_POSIT7346Output_9091);

SumNode_POSIT1745: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT7346Output_9091,ProductNode_POSIT7314Output_9053,SumNode_POSIT1745Output_9092);

ProductNode_POSIT7347: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1745Output_9092,ProductNode_POSIT7282Output_9015,ProductNode_POSIT7347Output_9093);

SumNode_POSIT1746: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT7347Output_9093,ProductNode_POSIT7243Output_8965,SumNode_POSIT1746Output_9094);

ProductNode_POSIT7348: entity work.PositMult_23_6_comb_uid2(arch)
port map(v13,SumNode_POSIT1746Output_9094,ProductNode_POSIT7348Output_9095);

ProductNode_POSIT7387: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1757Output_9144,ProductNode_POSIT6931Output_8579,ProductNode_POSIT7387Output_9145);

ProductNode_POSIT7414: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT7414weight,ProductNode_POSIT274Output_338,ProductNode_POSIT7414Output_9176);

ProductNode_POSIT7418: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT7418weight,ProductNode_POSIT278Output_343,ProductNode_POSIT7418Output_9181);

SumNode_POSIT1763: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT7418Output_9181,ProductNode_POSIT7414Output_9176,SumNode_POSIT1763Output_9182);

ProductNode_POSIT7419: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1763Output_9182,ProductNode_POSIT7201Output_8913,ProductNode_POSIT7419Output_9183);

ProductNode_POSIT7446: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT7446weight,ProductNode_POSIT274Output_338,ProductNode_POSIT7446Output_9214);

ProductNode_POSIT7450: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT7450weight,ProductNode_POSIT278Output_343,ProductNode_POSIT7450Output_9219);

SumNode_POSIT1769: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT7450Output_9219,ProductNode_POSIT7446Output_9214,SumNode_POSIT1769Output_9220);

ProductNode_POSIT7451: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1769Output_9220,ProductNode_POSIT7233Output_8951,ProductNode_POSIT7451Output_9221);

SumNode_POSIT1770: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT7451Output_9221,ProductNode_POSIT7419Output_9183,SumNode_POSIT1770Output_9222);

ProductNode_POSIT7452: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1770Output_9222,ProductNode_POSIT7387Output_9145,ProductNode_POSIT7452Output_9223);

ProductNode_POSIT7491: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1781Output_9272,ProductNode_POSIT7035Output_8707,ProductNode_POSIT7491Output_9273);

ProductNode_POSIT7518: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT7518weight,ProductNode_POSIT274Output_338,ProductNode_POSIT7518Output_9304);

ProductNode_POSIT7522: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT7522weight,ProductNode_POSIT278Output_343,ProductNode_POSIT7522Output_9309);

SumNode_POSIT1787: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT7522Output_9309,ProductNode_POSIT7518Output_9304,SumNode_POSIT1787Output_9310);

ProductNode_POSIT7523: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1787Output_9310,ProductNode_POSIT7305Output_9041,ProductNode_POSIT7523Output_9311);

ProductNode_POSIT7550: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT7550weight,ProductNode_POSIT274Output_338,ProductNode_POSIT7550Output_9342);

ProductNode_POSIT7554: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT7554weight,ProductNode_POSIT278Output_343,ProductNode_POSIT7554Output_9347);

SumNode_POSIT1793: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT7554Output_9347,ProductNode_POSIT7550Output_9342,SumNode_POSIT1793Output_9348);

ProductNode_POSIT7555: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1793Output_9348,ProductNode_POSIT7337Output_9079,ProductNode_POSIT7555Output_9349);

SumNode_POSIT1794: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT7555Output_9349,ProductNode_POSIT7523Output_9311,SumNode_POSIT1794Output_9350);

ProductNode_POSIT7556: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1794Output_9350,ProductNode_POSIT7491Output_9273,ProductNode_POSIT7556Output_9351);

SumNode_POSIT1795: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT7556Output_9351,ProductNode_POSIT7452Output_9223,SumNode_POSIT1795Output_9352);

ProductNode_POSIT7557: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb13,SumNode_POSIT1795Output_9352,ProductNode_POSIT7557Output_9353);

SumNode_POSIT1796: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT7557Output_9353,ProductNode_POSIT7348Output_9095,SumNode_POSIT1796Output_9354);

ProductNode_POSIT7558: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb3,SumNode_POSIT1796Output_9354,ProductNode_POSIT7558Output_9355);

SumNode_POSIT1797: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT7558Output_9355,ProductNode_POSIT7139Output_8837,SumNode_POSIT1797Output_9356);

ProductNode_POSIT7559: entity work.PositMult_23_6_comb_uid2(arch)
port map(v4,SumNode_POSIT1797Output_9356,ProductNode_POSIT7559Output_9357);

ProductNode_POSIT7561: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT7561weight,ProductNode_POSIT840Output_1039,ProductNode_POSIT7561Output_9359);

ProductNode_POSIT7570: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1799Output_9369,ProductNode_POSIT845Output_1045,ProductNode_POSIT7570Output_9370);

ProductNode_POSIT7578: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1801Output_9379,ProductNode_POSIT853Output_1055,ProductNode_POSIT7578Output_9380);

SumNode_POSIT1802: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT7578Output_9380,ProductNode_POSIT7570Output_9370,SumNode_POSIT1802Output_9381);

ProductNode_POSIT7579: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1802Output_9381,ProductNode_POSIT842Output_1041,ProductNode_POSIT7579Output_9382);

ProductNode_POSIT7588: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1804Output_9392,ProductNode_POSIT845Output_1045,ProductNode_POSIT7588Output_9393);

ProductNode_POSIT7596: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1806Output_9402,ProductNode_POSIT853Output_1055,ProductNode_POSIT7596Output_9403);

SumNode_POSIT1807: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT7596Output_9403,ProductNode_POSIT7588Output_9393,SumNode_POSIT1807Output_9404);

ProductNode_POSIT7597: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1807Output_9404,ProductNode_POSIT860Output_1064,ProductNode_POSIT7597Output_9405);

SumNode_POSIT1808: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT7597Output_9405,ProductNode_POSIT7579Output_9382,SumNode_POSIT1808Output_9406);

ProductNode_POSIT7598: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1808Output_9406,ProductNode_POSIT7561Output_9359,ProductNode_POSIT7598Output_9407);

ProductNode_POSIT7620: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT212Output_1112,ProductNode_POSIT6760Output_8370,ProductNode_POSIT7620Output_9432);

ProductNode_POSIT7621: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT7621weight,ProductNode_POSIT7620Output_9432,ProductNode_POSIT7621Output_9433);

ProductNode_POSIT7625: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT7625weight,ProductNode_POSIT904Output_1118,ProductNode_POSIT7625Output_9438);

ProductNode_POSIT7629: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT7629weight,ProductNode_POSIT908Output_1123,ProductNode_POSIT7629Output_9443);

SumNode_POSIT1814: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT7629Output_9443,ProductNode_POSIT7625Output_9438,SumNode_POSIT1814Output_9444);

ProductNode_POSIT7630: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1814Output_9444,ProductNode_POSIT7621Output_9433,ProductNode_POSIT7630Output_9445);

ProductNode_POSIT7652: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT218Output_1150,ProductNode_POSIT6792Output_8408,ProductNode_POSIT7652Output_9470);

ProductNode_POSIT7653: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT7653weight,ProductNode_POSIT7652Output_9470,ProductNode_POSIT7653Output_9471);

ProductNode_POSIT7657: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT7657weight,ProductNode_POSIT904Output_1118,ProductNode_POSIT7657Output_9476);

ProductNode_POSIT7661: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT7661weight,ProductNode_POSIT908Output_1123,ProductNode_POSIT7661Output_9481);

SumNode_POSIT1820: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT7661Output_9481,ProductNode_POSIT7657Output_9476,SumNode_POSIT1820Output_9482);

ProductNode_POSIT7662: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1820Output_9482,ProductNode_POSIT7653Output_9471,ProductNode_POSIT7662Output_9483);

SumNode_POSIT1821: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT7662Output_9483,ProductNode_POSIT7630Output_9445,SumNode_POSIT1821Output_9484);

ProductNode_POSIT7663: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1821Output_9484,ProductNode_POSIT7598Output_9407,ProductNode_POSIT7663Output_9485);

ProductNode_POSIT7665: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT7665weight,ProductNode_POSIT944Output_1167,ProductNode_POSIT7665Output_9487);

ProductNode_POSIT7674: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1823Output_9497,ProductNode_POSIT845Output_1045,ProductNode_POSIT7674Output_9498);

ProductNode_POSIT7682: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1825Output_9507,ProductNode_POSIT853Output_1055,ProductNode_POSIT7682Output_9508);

SumNode_POSIT1826: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT7682Output_9508,ProductNode_POSIT7674Output_9498,SumNode_POSIT1826Output_9509);

ProductNode_POSIT7683: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1826Output_9509,ProductNode_POSIT842Output_1041,ProductNode_POSIT7683Output_9510);

ProductNode_POSIT7692: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1828Output_9520,ProductNode_POSIT845Output_1045,ProductNode_POSIT7692Output_9521);

ProductNode_POSIT7700: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1830Output_9530,ProductNode_POSIT853Output_1055,ProductNode_POSIT7700Output_9531);

SumNode_POSIT1831: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT7700Output_9531,ProductNode_POSIT7692Output_9521,SumNode_POSIT1831Output_9532);

ProductNode_POSIT7701: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1831Output_9532,ProductNode_POSIT860Output_1064,ProductNode_POSIT7701Output_9533);

SumNode_POSIT1832: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT7701Output_9533,ProductNode_POSIT7683Output_9510,SumNode_POSIT1832Output_9534);

ProductNode_POSIT7702: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1832Output_9534,ProductNode_POSIT7665Output_9487,ProductNode_POSIT7702Output_9535);

ProductNode_POSIT7725: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT7725weight,ProductNode_POSIT7620Output_9432,ProductNode_POSIT7725Output_9561);

ProductNode_POSIT7729: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT7729weight,ProductNode_POSIT904Output_1118,ProductNode_POSIT7729Output_9566);

ProductNode_POSIT7733: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT7733weight,ProductNode_POSIT908Output_1123,ProductNode_POSIT7733Output_9571);

SumNode_POSIT1838: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT7733Output_9571,ProductNode_POSIT7729Output_9566,SumNode_POSIT1838Output_9572);

ProductNode_POSIT7734: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1838Output_9572,ProductNode_POSIT7725Output_9561,ProductNode_POSIT7734Output_9573);

ProductNode_POSIT7757: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT7757weight,ProductNode_POSIT7652Output_9470,ProductNode_POSIT7757Output_9599);

ProductNode_POSIT7761: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT7761weight,ProductNode_POSIT904Output_1118,ProductNode_POSIT7761Output_9604);

ProductNode_POSIT7765: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT7765weight,ProductNode_POSIT908Output_1123,ProductNode_POSIT7765Output_9609);

SumNode_POSIT1844: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT7765Output_9609,ProductNode_POSIT7761Output_9604,SumNode_POSIT1844Output_9610);

ProductNode_POSIT7766: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1844Output_9610,ProductNode_POSIT7757Output_9599,ProductNode_POSIT7766Output_9611);

SumNode_POSIT1845: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT7766Output_9611,ProductNode_POSIT7734Output_9573,SumNode_POSIT1845Output_9612);

ProductNode_POSIT7767: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1845Output_9612,ProductNode_POSIT7702Output_9535,ProductNode_POSIT7767Output_9613);

SumNode_POSIT1846: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT7767Output_9613,ProductNode_POSIT7663Output_9485,SumNode_POSIT1846Output_9614);

ProductNode_POSIT7768: entity work.PositMult_23_6_comb_uid2(arch)
port map(v13,SumNode_POSIT1846Output_9614,ProductNode_POSIT7768Output_9615);

ProductNode_POSIT7770: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT7770weight,ProductNode_POSIT840Output_1039,ProductNode_POSIT7770Output_9617);

ProductNode_POSIT7807: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1857Output_9664,ProductNode_POSIT7770Output_9617,ProductNode_POSIT7807Output_9665);

ProductNode_POSIT7834: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT7834weight,ProductNode_POSIT1113Output_1376,ProductNode_POSIT7834Output_9696);

ProductNode_POSIT7838: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT7838weight,ProductNode_POSIT1117Output_1381,ProductNode_POSIT7838Output_9701);

SumNode_POSIT1863: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT7838Output_9701,ProductNode_POSIT7834Output_9696,SumNode_POSIT1863Output_9702);

ProductNode_POSIT7839: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1863Output_9702,ProductNode_POSIT7621Output_9433,ProductNode_POSIT7839Output_9703);

ProductNode_POSIT7866: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT7866weight,ProductNode_POSIT1113Output_1376,ProductNode_POSIT7866Output_9734);

ProductNode_POSIT7870: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT7870weight,ProductNode_POSIT1117Output_1381,ProductNode_POSIT7870Output_9739);

SumNode_POSIT1869: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT7870Output_9739,ProductNode_POSIT7866Output_9734,SumNode_POSIT1869Output_9740);

ProductNode_POSIT7871: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1869Output_9740,ProductNode_POSIT7653Output_9471,ProductNode_POSIT7871Output_9741);

SumNode_POSIT1870: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT7871Output_9741,ProductNode_POSIT7839Output_9703,SumNode_POSIT1870Output_9742);

ProductNode_POSIT7872: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1870Output_9742,ProductNode_POSIT7807Output_9665,ProductNode_POSIT7872Output_9743);

ProductNode_POSIT7874: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT7874weight,ProductNode_POSIT944Output_1167,ProductNode_POSIT7874Output_9745);

ProductNode_POSIT7911: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1881Output_9792,ProductNode_POSIT7874Output_9745,ProductNode_POSIT7911Output_9793);

ProductNode_POSIT7938: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT7938weight,ProductNode_POSIT1113Output_1376,ProductNode_POSIT7938Output_9824);

ProductNode_POSIT7942: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT7942weight,ProductNode_POSIT1117Output_1381,ProductNode_POSIT7942Output_9829);

SumNode_POSIT1887: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT7942Output_9829,ProductNode_POSIT7938Output_9824,SumNode_POSIT1887Output_9830);

ProductNode_POSIT7943: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1887Output_9830,ProductNode_POSIT7725Output_9561,ProductNode_POSIT7943Output_9831);

ProductNode_POSIT7970: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT7970weight,ProductNode_POSIT1113Output_1376,ProductNode_POSIT7970Output_9862);

ProductNode_POSIT7974: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT7974weight,ProductNode_POSIT1117Output_1381,ProductNode_POSIT7974Output_9867);

SumNode_POSIT1893: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT7974Output_9867,ProductNode_POSIT7970Output_9862,SumNode_POSIT1893Output_9868);

ProductNode_POSIT7975: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1893Output_9868,ProductNode_POSIT7757Output_9599,ProductNode_POSIT7975Output_9869);

SumNode_POSIT1894: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT7975Output_9869,ProductNode_POSIT7943Output_9831,SumNode_POSIT1894Output_9870);

ProductNode_POSIT7976: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1894Output_9870,ProductNode_POSIT7911Output_9793,ProductNode_POSIT7976Output_9871);

SumNode_POSIT1895: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT7976Output_9871,ProductNode_POSIT7872Output_9743,SumNode_POSIT1895Output_9872);

ProductNode_POSIT7977: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb13,SumNode_POSIT1895Output_9872,ProductNode_POSIT7977Output_9873);

SumNode_POSIT1896: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT7977Output_9873,ProductNode_POSIT7768Output_9615,SumNode_POSIT1896Output_9874);

ProductNode_POSIT7978: entity work.PositMult_23_6_comb_uid2(arch)
port map(v3,SumNode_POSIT1896Output_9874,ProductNode_POSIT7978Output_9875);

ProductNode_POSIT7998: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1901Output_9899,ProductNode_POSIT1261Output_1559,ProductNode_POSIT7998Output_9900);

ProductNode_POSIT8016: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1906Output_9922,ProductNode_POSIT1279Output_1582,ProductNode_POSIT8016Output_9923);

SumNode_POSIT1907: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT8016Output_9923,ProductNode_POSIT7998Output_9900,SumNode_POSIT1907Output_9924);

ProductNode_POSIT8017: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1907Output_9924,ProductNode_POSIT7561Output_9359,ProductNode_POSIT8017Output_9925);

ProductNode_POSIT8039: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT311Output_1630,ProductNode_POSIT6760Output_8370,ProductNode_POSIT8039Output_9950);

ProductNode_POSIT8040: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT8040weight,ProductNode_POSIT8039Output_9950,ProductNode_POSIT8040Output_9951);

ProductNode_POSIT8044: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT8044weight,ProductNode_POSIT904Output_1118,ProductNode_POSIT8044Output_9956);

ProductNode_POSIT8048: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT8048weight,ProductNode_POSIT908Output_1123,ProductNode_POSIT8048Output_9961);

SumNode_POSIT1913: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT8048Output_9961,ProductNode_POSIT8044Output_9956,SumNode_POSIT1913Output_9962);

ProductNode_POSIT8049: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1913Output_9962,ProductNode_POSIT8040Output_9951,ProductNode_POSIT8049Output_9963);

ProductNode_POSIT8071: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT317Output_1668,ProductNode_POSIT6792Output_8408,ProductNode_POSIT8071Output_9988);

ProductNode_POSIT8072: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT8072weight,ProductNode_POSIT8071Output_9988,ProductNode_POSIT8072Output_9989);

ProductNode_POSIT8076: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT8076weight,ProductNode_POSIT904Output_1118,ProductNode_POSIT8076Output_9994);

ProductNode_POSIT8080: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT8080weight,ProductNode_POSIT908Output_1123,ProductNode_POSIT8080Output_9999);

SumNode_POSIT1919: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT8080Output_9999,ProductNode_POSIT8076Output_9994,SumNode_POSIT1919Output_10000);

ProductNode_POSIT8081: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1919Output_10000,ProductNode_POSIT8072Output_9989,ProductNode_POSIT8081Output_10001);

SumNode_POSIT1920: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT8081Output_10001,ProductNode_POSIT8049Output_9963,SumNode_POSIT1920Output_10002);

ProductNode_POSIT8082: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1920Output_10002,ProductNode_POSIT8017Output_9925,ProductNode_POSIT8082Output_10003);

ProductNode_POSIT8102: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1925Output_10027,ProductNode_POSIT1261Output_1559,ProductNode_POSIT8102Output_10028);

ProductNode_POSIT8120: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1930Output_10050,ProductNode_POSIT1279Output_1582,ProductNode_POSIT8120Output_10051);

SumNode_POSIT1931: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT8120Output_10051,ProductNode_POSIT8102Output_10028,SumNode_POSIT1931Output_10052);

ProductNode_POSIT8121: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1931Output_10052,ProductNode_POSIT7665Output_9487,ProductNode_POSIT8121Output_10053);

ProductNode_POSIT8144: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT8144weight,ProductNode_POSIT8039Output_9950,ProductNode_POSIT8144Output_10079);

ProductNode_POSIT8148: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT8148weight,ProductNode_POSIT904Output_1118,ProductNode_POSIT8148Output_10084);

ProductNode_POSIT8152: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT8152weight,ProductNode_POSIT908Output_1123,ProductNode_POSIT8152Output_10089);

SumNode_POSIT1937: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT8152Output_10089,ProductNode_POSIT8148Output_10084,SumNode_POSIT1937Output_10090);

ProductNode_POSIT8153: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1937Output_10090,ProductNode_POSIT8144Output_10079,ProductNode_POSIT8153Output_10091);

ProductNode_POSIT8176: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT8176weight,ProductNode_POSIT8071Output_9988,ProductNode_POSIT8176Output_10117);

ProductNode_POSIT8180: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT8180weight,ProductNode_POSIT904Output_1118,ProductNode_POSIT8180Output_10122);

ProductNode_POSIT8184: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT8184weight,ProductNode_POSIT908Output_1123,ProductNode_POSIT8184Output_10127);

SumNode_POSIT1943: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT8184Output_10127,ProductNode_POSIT8180Output_10122,SumNode_POSIT1943Output_10128);

ProductNode_POSIT8185: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1943Output_10128,ProductNode_POSIT8176Output_10117,ProductNode_POSIT8185Output_10129);

SumNode_POSIT1944: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT8185Output_10129,ProductNode_POSIT8153Output_10091,SumNode_POSIT1944Output_10130);

ProductNode_POSIT8186: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1944Output_10130,ProductNode_POSIT8121Output_10053,ProductNode_POSIT8186Output_10131);

SumNode_POSIT1945: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT8186Output_10131,ProductNode_POSIT8082Output_10003,SumNode_POSIT1945Output_10132);

ProductNode_POSIT8187: entity work.PositMult_23_6_comb_uid2(arch)
port map(v13,SumNode_POSIT1945Output_10132,ProductNode_POSIT8187Output_10133);

ProductNode_POSIT8226: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1956Output_10182,ProductNode_POSIT7770Output_9617,ProductNode_POSIT8226Output_10183);

ProductNode_POSIT8253: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT8253weight,ProductNode_POSIT1113Output_1376,ProductNode_POSIT8253Output_10214);

ProductNode_POSIT8257: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT8257weight,ProductNode_POSIT1117Output_1381,ProductNode_POSIT8257Output_10219);

SumNode_POSIT1962: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT8257Output_10219,ProductNode_POSIT8253Output_10214,SumNode_POSIT1962Output_10220);

ProductNode_POSIT8258: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1962Output_10220,ProductNode_POSIT8040Output_9951,ProductNode_POSIT8258Output_10221);

ProductNode_POSIT8285: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT8285weight,ProductNode_POSIT1113Output_1376,ProductNode_POSIT8285Output_10252);

ProductNode_POSIT8289: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT8289weight,ProductNode_POSIT1117Output_1381,ProductNode_POSIT8289Output_10257);

SumNode_POSIT1968: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT8289Output_10257,ProductNode_POSIT8285Output_10252,SumNode_POSIT1968Output_10258);

ProductNode_POSIT8290: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1968Output_10258,ProductNode_POSIT8072Output_9989,ProductNode_POSIT8290Output_10259);

SumNode_POSIT1969: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT8290Output_10259,ProductNode_POSIT8258Output_10221,SumNode_POSIT1969Output_10260);

ProductNode_POSIT8291: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1969Output_10260,ProductNode_POSIT8226Output_10183,ProductNode_POSIT8291Output_10261);

ProductNode_POSIT8330: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1980Output_10310,ProductNode_POSIT7874Output_9745,ProductNode_POSIT8330Output_10311);

ProductNode_POSIT8357: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT8357weight,ProductNode_POSIT1113Output_1376,ProductNode_POSIT8357Output_10342);

ProductNode_POSIT8361: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT8361weight,ProductNode_POSIT1117Output_1381,ProductNode_POSIT8361Output_10347);

SumNode_POSIT1986: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT8361Output_10347,ProductNode_POSIT8357Output_10342,SumNode_POSIT1986Output_10348);

ProductNode_POSIT8362: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1986Output_10348,ProductNode_POSIT8144Output_10079,ProductNode_POSIT8362Output_10349);

ProductNode_POSIT8389: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT8389weight,ProductNode_POSIT1113Output_1376,ProductNode_POSIT8389Output_10380);

ProductNode_POSIT8393: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT8393weight,ProductNode_POSIT1117Output_1381,ProductNode_POSIT8393Output_10385);

SumNode_POSIT1992: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT8393Output_10385,ProductNode_POSIT8389Output_10380,SumNode_POSIT1992Output_10386);

ProductNode_POSIT8394: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1992Output_10386,ProductNode_POSIT8176Output_10117,ProductNode_POSIT8394Output_10387);

SumNode_POSIT1993: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT8394Output_10387,ProductNode_POSIT8362Output_10349,SumNode_POSIT1993Output_10388);

ProductNode_POSIT8395: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1993Output_10388,ProductNode_POSIT8330Output_10311,ProductNode_POSIT8395Output_10389);

SumNode_POSIT1994: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT8395Output_10389,ProductNode_POSIT8291Output_10261,SumNode_POSIT1994Output_10390);

ProductNode_POSIT8396: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb13,SumNode_POSIT1994Output_10390,ProductNode_POSIT8396Output_10391);

SumNode_POSIT1995: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT8396Output_10391,ProductNode_POSIT8187Output_10133,SumNode_POSIT1995Output_10392);

ProductNode_POSIT8397: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb3,SumNode_POSIT1995Output_10392,ProductNode_POSIT8397Output_10393);

SumNode_POSIT1996: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT8397Output_10393,ProductNode_POSIT7978Output_9875,SumNode_POSIT1996Output_10394);

ProductNode_POSIT8398: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb4,SumNode_POSIT1996Output_10394,ProductNode_POSIT8398Output_10395);

SumNode_POSIT1997: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT8398Output_10395,ProductNode_POSIT7559Output_9357,SumNode_POSIT1997Output_10396);

ProductNode_POSIT8399: entity work.PositMult_23_6_comb_uid2(arch)
port map(v12,SumNode_POSIT1997Output_10396,ProductNode_POSIT8399Output_10397);

ProductNode_POSIT8401: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT8401weight,ProductNode_POSIT1680Output_2079,ProductNode_POSIT8401Output_10399);

ProductNode_POSIT8407: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT8407weight,ProductNode_POSIT1686Output_2086,ProductNode_POSIT8407Output_10406);

ProductNode_POSIT8409: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT8409weight,ProductNode_POSIT1688Output_2088,ProductNode_POSIT8409Output_10408);

SumNode_POSIT1999: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT8409Output_10408,ProductNode_POSIT8407Output_10406,SumNode_POSIT1999Output_10409);

ProductNode_POSIT8410: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1999Output_10409,ProductNode_POSIT1685Output_2085,ProductNode_POSIT8410Output_10410);

ProductNode_POSIT8415: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT8415weight,ProductNode_POSIT1694Output_2096,ProductNode_POSIT8415Output_10416);

ProductNode_POSIT8417: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT8417weight,ProductNode_POSIT1696Output_2098,ProductNode_POSIT8417Output_10418);

SumNode_POSIT2001: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT8417Output_10418,ProductNode_POSIT8415Output_10416,SumNode_POSIT2001Output_10419);

ProductNode_POSIT8418: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2001Output_10419,ProductNode_POSIT1693Output_2095,ProductNode_POSIT8418Output_10420);

SumNode_POSIT2002: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT8418Output_10420,ProductNode_POSIT8410Output_10410,SumNode_POSIT2002Output_10421);

ProductNode_POSIT8419: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2002Output_10421,ProductNode_POSIT1682Output_2081,ProductNode_POSIT8419Output_10422);

ProductNode_POSIT8425: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT8425weight,ProductNode_POSIT1704Output_2109,ProductNode_POSIT8425Output_10429);

ProductNode_POSIT8427: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT8427weight,ProductNode_POSIT1706Output_2111,ProductNode_POSIT8427Output_10431);

SumNode_POSIT2004: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT8427Output_10431,ProductNode_POSIT8425Output_10429,SumNode_POSIT2004Output_10432);

ProductNode_POSIT8428: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2004Output_10432,ProductNode_POSIT1685Output_2085,ProductNode_POSIT8428Output_10433);

ProductNode_POSIT8433: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT8433weight,ProductNode_POSIT1712Output_2119,ProductNode_POSIT8433Output_10439);

ProductNode_POSIT8435: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT8435weight,ProductNode_POSIT1714Output_2121,ProductNode_POSIT8435Output_10441);

SumNode_POSIT2006: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT8435Output_10441,ProductNode_POSIT8433Output_10439,SumNode_POSIT2006Output_10442);

ProductNode_POSIT8436: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2006Output_10442,ProductNode_POSIT1693Output_2095,ProductNode_POSIT8436Output_10443);

SumNode_POSIT2007: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT8436Output_10443,ProductNode_POSIT8428Output_10433,SumNode_POSIT2007Output_10444);

ProductNode_POSIT8437: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2007Output_10444,ProductNode_POSIT1700Output_2104,ProductNode_POSIT8437Output_10445);

SumNode_POSIT2008: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT8437Output_10445,ProductNode_POSIT8419Output_10422,SumNode_POSIT2008Output_10446);

ProductNode_POSIT8438: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2008Output_10446,ProductNode_POSIT8401Output_10399,ProductNode_POSIT8438Output_10447);

ProductNode_POSIT8465: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT8465weight,ProductNode_POSIT1744Output_2158,ProductNode_POSIT8465Output_10478);

ProductNode_POSIT8469: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT8469weight,ProductNode_POSIT278Output_343,ProductNode_POSIT8469Output_10483);

SumNode_POSIT2014: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT8469Output_10483,ProductNode_POSIT8465Output_10478,SumNode_POSIT2014Output_10484);

ProductNode_POSIT8470: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2014Output_10484,ProductNode_POSIT6782Output_8395,ProductNode_POSIT8470Output_10485);

ProductNode_POSIT8497: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT8497weight,ProductNode_POSIT1744Output_2158,ProductNode_POSIT8497Output_10516);

ProductNode_POSIT8501: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT8501weight,ProductNode_POSIT278Output_343,ProductNode_POSIT8501Output_10521);

SumNode_POSIT2020: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT8501Output_10521,ProductNode_POSIT8497Output_10516,SumNode_POSIT2020Output_10522);

ProductNode_POSIT8502: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2020Output_10522,ProductNode_POSIT6814Output_8433,ProductNode_POSIT8502Output_10523);

SumNode_POSIT2021: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT8502Output_10523,ProductNode_POSIT8470Output_10485,SumNode_POSIT2021Output_10524);

ProductNode_POSIT8503: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2021Output_10524,ProductNode_POSIT8438Output_10447,ProductNode_POSIT8503Output_10525);

ProductNode_POSIT8505: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT8505weight,ProductNode_POSIT1784Output_2207,ProductNode_POSIT8505Output_10527);

ProductNode_POSIT8511: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT8511weight,ProductNode_POSIT1686Output_2086,ProductNode_POSIT8511Output_10534);

ProductNode_POSIT8513: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT8513weight,ProductNode_POSIT1688Output_2088,ProductNode_POSIT8513Output_10536);

SumNode_POSIT2023: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT8513Output_10536,ProductNode_POSIT8511Output_10534,SumNode_POSIT2023Output_10537);

ProductNode_POSIT8514: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2023Output_10537,ProductNode_POSIT1685Output_2085,ProductNode_POSIT8514Output_10538);

ProductNode_POSIT8519: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT8519weight,ProductNode_POSIT1694Output_2096,ProductNode_POSIT8519Output_10544);

ProductNode_POSIT8521: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT8521weight,ProductNode_POSIT1696Output_2098,ProductNode_POSIT8521Output_10546);

SumNode_POSIT2025: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT8521Output_10546,ProductNode_POSIT8519Output_10544,SumNode_POSIT2025Output_10547);

ProductNode_POSIT8522: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2025Output_10547,ProductNode_POSIT1693Output_2095,ProductNode_POSIT8522Output_10548);

SumNode_POSIT2026: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT8522Output_10548,ProductNode_POSIT8514Output_10538,SumNode_POSIT2026Output_10549);

ProductNode_POSIT8523: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2026Output_10549,ProductNode_POSIT1682Output_2081,ProductNode_POSIT8523Output_10550);

ProductNode_POSIT8529: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT8529weight,ProductNode_POSIT1704Output_2109,ProductNode_POSIT8529Output_10557);

ProductNode_POSIT8531: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT8531weight,ProductNode_POSIT1706Output_2111,ProductNode_POSIT8531Output_10559);

SumNode_POSIT2028: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT8531Output_10559,ProductNode_POSIT8529Output_10557,SumNode_POSIT2028Output_10560);

ProductNode_POSIT8532: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2028Output_10560,ProductNode_POSIT1685Output_2085,ProductNode_POSIT8532Output_10561);

ProductNode_POSIT8537: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT8537weight,ProductNode_POSIT1712Output_2119,ProductNode_POSIT8537Output_10567);

ProductNode_POSIT8539: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT8539weight,ProductNode_POSIT1714Output_2121,ProductNode_POSIT8539Output_10569);

SumNode_POSIT2030: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT8539Output_10569,ProductNode_POSIT8537Output_10567,SumNode_POSIT2030Output_10570);

ProductNode_POSIT8540: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2030Output_10570,ProductNode_POSIT1693Output_2095,ProductNode_POSIT8540Output_10571);

SumNode_POSIT2031: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT8540Output_10571,ProductNode_POSIT8532Output_10561,SumNode_POSIT2031Output_10572);

ProductNode_POSIT8541: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2031Output_10572,ProductNode_POSIT1700Output_2104,ProductNode_POSIT8541Output_10573);

SumNode_POSIT2032: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT8541Output_10573,ProductNode_POSIT8523Output_10550,SumNode_POSIT2032Output_10574);

ProductNode_POSIT8542: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2032Output_10574,ProductNode_POSIT8505Output_10527,ProductNode_POSIT8542Output_10575);

ProductNode_POSIT8569: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT8569weight,ProductNode_POSIT1744Output_2158,ProductNode_POSIT8569Output_10606);

ProductNode_POSIT8573: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT8573weight,ProductNode_POSIT278Output_343,ProductNode_POSIT8573Output_10611);

SumNode_POSIT2038: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT8573Output_10611,ProductNode_POSIT8569Output_10606,SumNode_POSIT2038Output_10612);

ProductNode_POSIT8574: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2038Output_10612,ProductNode_POSIT6886Output_8523,ProductNode_POSIT8574Output_10613);

ProductNode_POSIT8601: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT8601weight,ProductNode_POSIT1744Output_2158,ProductNode_POSIT8601Output_10644);

ProductNode_POSIT8605: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT8605weight,ProductNode_POSIT278Output_343,ProductNode_POSIT8605Output_10649);

SumNode_POSIT2044: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT8605Output_10649,ProductNode_POSIT8601Output_10644,SumNode_POSIT2044Output_10650);

ProductNode_POSIT8606: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2044Output_10650,ProductNode_POSIT6918Output_8561,ProductNode_POSIT8606Output_10651);

SumNode_POSIT2045: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT8606Output_10651,ProductNode_POSIT8574Output_10613,SumNode_POSIT2045Output_10652);

ProductNode_POSIT8607: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2045Output_10652,ProductNode_POSIT8542Output_10575,ProductNode_POSIT8607Output_10653);

SumNode_POSIT2046: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT8607Output_10653,ProductNode_POSIT8503Output_10525,SumNode_POSIT2046Output_10654);

ProductNode_POSIT8608: entity work.PositMult_23_6_comb_uid2(arch)
port map(v13,SumNode_POSIT2046Output_10654,ProductNode_POSIT8608Output_10655);

ProductNode_POSIT8610: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT8610weight,ProductNode_POSIT1680Output_2079,ProductNode_POSIT8610Output_10657);

ProductNode_POSIT8647: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2057Output_10704,ProductNode_POSIT8610Output_10657,ProductNode_POSIT8647Output_10705);

ProductNode_POSIT8674: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT8674weight,ProductNode_POSIT1953Output_2416,ProductNode_POSIT8674Output_10736);

ProductNode_POSIT8678: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT8678weight,ProductNode_POSIT1957Output_2421,ProductNode_POSIT8678Output_10741);

SumNode_POSIT2063: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT8678Output_10741,ProductNode_POSIT8674Output_10736,SumNode_POSIT2063Output_10742);

ProductNode_POSIT8679: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2063Output_10742,ProductNode_POSIT6782Output_8395,ProductNode_POSIT8679Output_10743);

ProductNode_POSIT8706: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT8706weight,ProductNode_POSIT1953Output_2416,ProductNode_POSIT8706Output_10774);

ProductNode_POSIT8710: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT8710weight,ProductNode_POSIT1957Output_2421,ProductNode_POSIT8710Output_10779);

SumNode_POSIT2069: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT8710Output_10779,ProductNode_POSIT8706Output_10774,SumNode_POSIT2069Output_10780);

ProductNode_POSIT8711: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2069Output_10780,ProductNode_POSIT6814Output_8433,ProductNode_POSIT8711Output_10781);

SumNode_POSIT2070: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT8711Output_10781,ProductNode_POSIT8679Output_10743,SumNode_POSIT2070Output_10782);

ProductNode_POSIT8712: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2070Output_10782,ProductNode_POSIT8647Output_10705,ProductNode_POSIT8712Output_10783);

ProductNode_POSIT8714: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT8714weight,ProductNode_POSIT1784Output_2207,ProductNode_POSIT8714Output_10785);

ProductNode_POSIT8751: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2081Output_10832,ProductNode_POSIT8714Output_10785,ProductNode_POSIT8751Output_10833);

ProductNode_POSIT8778: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT8778weight,ProductNode_POSIT1953Output_2416,ProductNode_POSIT8778Output_10864);

ProductNode_POSIT8782: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT8782weight,ProductNode_POSIT1957Output_2421,ProductNode_POSIT8782Output_10869);

SumNode_POSIT2087: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT8782Output_10869,ProductNode_POSIT8778Output_10864,SumNode_POSIT2087Output_10870);

ProductNode_POSIT8783: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2087Output_10870,ProductNode_POSIT6886Output_8523,ProductNode_POSIT8783Output_10871);

ProductNode_POSIT8810: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT8810weight,ProductNode_POSIT1953Output_2416,ProductNode_POSIT8810Output_10902);

ProductNode_POSIT8814: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT8814weight,ProductNode_POSIT1957Output_2421,ProductNode_POSIT8814Output_10907);

SumNode_POSIT2093: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT8814Output_10907,ProductNode_POSIT8810Output_10902,SumNode_POSIT2093Output_10908);

ProductNode_POSIT8815: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2093Output_10908,ProductNode_POSIT6918Output_8561,ProductNode_POSIT8815Output_10909);

SumNode_POSIT2094: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT8815Output_10909,ProductNode_POSIT8783Output_10871,SumNode_POSIT2094Output_10910);

ProductNode_POSIT8816: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2094Output_10910,ProductNode_POSIT8751Output_10833,ProductNode_POSIT8816Output_10911);

SumNode_POSIT2095: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT8816Output_10911,ProductNode_POSIT8712Output_10783,SumNode_POSIT2095Output_10912);

ProductNode_POSIT8817: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb13,SumNode_POSIT2095Output_10912,ProductNode_POSIT8817Output_10913);

SumNode_POSIT2096: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT8817Output_10913,ProductNode_POSIT8608Output_10655,SumNode_POSIT2096Output_10914);

ProductNode_POSIT8818: entity work.PositMult_23_6_comb_uid2(arch)
port map(v3,SumNode_POSIT2096Output_10914,ProductNode_POSIT8818Output_10915);

ProductNode_POSIT8838: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2101Output_10939,ProductNode_POSIT2101Output_2599,ProductNode_POSIT8838Output_10940);

ProductNode_POSIT8856: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2106Output_10962,ProductNode_POSIT2119Output_2622,ProductNode_POSIT8856Output_10963);

SumNode_POSIT2107: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT8856Output_10963,ProductNode_POSIT8838Output_10940,SumNode_POSIT2107Output_10964);

ProductNode_POSIT8857: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2107Output_10964,ProductNode_POSIT8401Output_10399,ProductNode_POSIT8857Output_10965);

ProductNode_POSIT8884: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT8884weight,ProductNode_POSIT1744Output_2158,ProductNode_POSIT8884Output_10996);

ProductNode_POSIT8888: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT8888weight,ProductNode_POSIT278Output_343,ProductNode_POSIT8888Output_11001);

SumNode_POSIT2113: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT8888Output_11001,ProductNode_POSIT8884Output_10996,SumNode_POSIT2113Output_11002);

ProductNode_POSIT8889: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2113Output_11002,ProductNode_POSIT7201Output_8913,ProductNode_POSIT8889Output_11003);

ProductNode_POSIT8916: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT8916weight,ProductNode_POSIT1744Output_2158,ProductNode_POSIT8916Output_11034);

ProductNode_POSIT8920: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT8920weight,ProductNode_POSIT278Output_343,ProductNode_POSIT8920Output_11039);

SumNode_POSIT2119: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT8920Output_11039,ProductNode_POSIT8916Output_11034,SumNode_POSIT2119Output_11040);

ProductNode_POSIT8921: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2119Output_11040,ProductNode_POSIT7233Output_8951,ProductNode_POSIT8921Output_11041);

SumNode_POSIT2120: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT8921Output_11041,ProductNode_POSIT8889Output_11003,SumNode_POSIT2120Output_11042);

ProductNode_POSIT8922: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2120Output_11042,ProductNode_POSIT8857Output_10965,ProductNode_POSIT8922Output_11043);

ProductNode_POSIT8942: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2125Output_11067,ProductNode_POSIT2101Output_2599,ProductNode_POSIT8942Output_11068);

ProductNode_POSIT8960: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2130Output_11090,ProductNode_POSIT2119Output_2622,ProductNode_POSIT8960Output_11091);

SumNode_POSIT2131: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT8960Output_11091,ProductNode_POSIT8942Output_11068,SumNode_POSIT2131Output_11092);

ProductNode_POSIT8961: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2131Output_11092,ProductNode_POSIT8505Output_10527,ProductNode_POSIT8961Output_11093);

ProductNode_POSIT8988: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT8988weight,ProductNode_POSIT1744Output_2158,ProductNode_POSIT8988Output_11124);

ProductNode_POSIT8992: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT8992weight,ProductNode_POSIT278Output_343,ProductNode_POSIT8992Output_11129);

SumNode_POSIT2137: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT8992Output_11129,ProductNode_POSIT8988Output_11124,SumNode_POSIT2137Output_11130);

ProductNode_POSIT8993: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2137Output_11130,ProductNode_POSIT7305Output_9041,ProductNode_POSIT8993Output_11131);

ProductNode_POSIT9020: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT9020weight,ProductNode_POSIT1744Output_2158,ProductNode_POSIT9020Output_11162);

ProductNode_POSIT9024: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT9024weight,ProductNode_POSIT278Output_343,ProductNode_POSIT9024Output_11167);

SumNode_POSIT2143: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT9024Output_11167,ProductNode_POSIT9020Output_11162,SumNode_POSIT2143Output_11168);

ProductNode_POSIT9025: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2143Output_11168,ProductNode_POSIT7337Output_9079,ProductNode_POSIT9025Output_11169);

SumNode_POSIT2144: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT9025Output_11169,ProductNode_POSIT8993Output_11131,SumNode_POSIT2144Output_11170);

ProductNode_POSIT9026: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2144Output_11170,ProductNode_POSIT8961Output_11093,ProductNode_POSIT9026Output_11171);

SumNode_POSIT2145: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT9026Output_11171,ProductNode_POSIT8922Output_11043,SumNode_POSIT2145Output_11172);

ProductNode_POSIT9027: entity work.PositMult_23_6_comb_uid2(arch)
port map(v13,SumNode_POSIT2145Output_11172,ProductNode_POSIT9027Output_11173);

ProductNode_POSIT9066: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2156Output_11222,ProductNode_POSIT8610Output_10657,ProductNode_POSIT9066Output_11223);

ProductNode_POSIT9093: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT9093weight,ProductNode_POSIT1953Output_2416,ProductNode_POSIT9093Output_11254);

ProductNode_POSIT9097: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT9097weight,ProductNode_POSIT1957Output_2421,ProductNode_POSIT9097Output_11259);

SumNode_POSIT2162: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT9097Output_11259,ProductNode_POSIT9093Output_11254,SumNode_POSIT2162Output_11260);

ProductNode_POSIT9098: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2162Output_11260,ProductNode_POSIT7201Output_8913,ProductNode_POSIT9098Output_11261);

ProductNode_POSIT9125: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT9125weight,ProductNode_POSIT1953Output_2416,ProductNode_POSIT9125Output_11292);

ProductNode_POSIT9129: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT9129weight,ProductNode_POSIT1957Output_2421,ProductNode_POSIT9129Output_11297);

SumNode_POSIT2168: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT9129Output_11297,ProductNode_POSIT9125Output_11292,SumNode_POSIT2168Output_11298);

ProductNode_POSIT9130: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2168Output_11298,ProductNode_POSIT7233Output_8951,ProductNode_POSIT9130Output_11299);

SumNode_POSIT2169: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT9130Output_11299,ProductNode_POSIT9098Output_11261,SumNode_POSIT2169Output_11300);

ProductNode_POSIT9131: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2169Output_11300,ProductNode_POSIT9066Output_11223,ProductNode_POSIT9131Output_11301);

ProductNode_POSIT9170: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2180Output_11350,ProductNode_POSIT8714Output_10785,ProductNode_POSIT9170Output_11351);

ProductNode_POSIT9197: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT9197weight,ProductNode_POSIT1953Output_2416,ProductNode_POSIT9197Output_11382);

ProductNode_POSIT9201: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT9201weight,ProductNode_POSIT1957Output_2421,ProductNode_POSIT9201Output_11387);

SumNode_POSIT2186: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT9201Output_11387,ProductNode_POSIT9197Output_11382,SumNode_POSIT2186Output_11388);

ProductNode_POSIT9202: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2186Output_11388,ProductNode_POSIT7305Output_9041,ProductNode_POSIT9202Output_11389);

ProductNode_POSIT9229: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT9229weight,ProductNode_POSIT1953Output_2416,ProductNode_POSIT9229Output_11420);

ProductNode_POSIT9233: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT9233weight,ProductNode_POSIT1957Output_2421,ProductNode_POSIT9233Output_11425);

SumNode_POSIT2192: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT9233Output_11425,ProductNode_POSIT9229Output_11420,SumNode_POSIT2192Output_11426);

ProductNode_POSIT9234: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2192Output_11426,ProductNode_POSIT7337Output_9079,ProductNode_POSIT9234Output_11427);

SumNode_POSIT2193: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT9234Output_11427,ProductNode_POSIT9202Output_11389,SumNode_POSIT2193Output_11428);

ProductNode_POSIT9235: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2193Output_11428,ProductNode_POSIT9170Output_11351,ProductNode_POSIT9235Output_11429);

SumNode_POSIT2194: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT9235Output_11429,ProductNode_POSIT9131Output_11301,SumNode_POSIT2194Output_11430);

ProductNode_POSIT9236: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb13,SumNode_POSIT2194Output_11430,ProductNode_POSIT9236Output_11431);

SumNode_POSIT2195: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT9236Output_11431,ProductNode_POSIT9027Output_11173,SumNode_POSIT2195Output_11432);

ProductNode_POSIT9237: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb3,SumNode_POSIT2195Output_11432,ProductNode_POSIT9237Output_11433);

SumNode_POSIT2196: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT9237Output_11433,ProductNode_POSIT8818Output_10915,SumNode_POSIT2196Output_11434);

ProductNode_POSIT9238: entity work.PositMult_23_6_comb_uid2(arch)
port map(v4,SumNode_POSIT2196Output_11434,ProductNode_POSIT9238Output_11435);

ProductNode_POSIT9240: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT9240weight,ProductNode_POSIT2519Output_3117,ProductNode_POSIT9240Output_11437);

ProductNode_POSIT9249: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2198Output_11447,ProductNode_POSIT2524Output_3123,ProductNode_POSIT9249Output_11448);

ProductNode_POSIT9257: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2200Output_11457,ProductNode_POSIT2532Output_3133,ProductNode_POSIT9257Output_11458);

SumNode_POSIT2201: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT9257Output_11458,ProductNode_POSIT9249Output_11448,SumNode_POSIT2201Output_11459);

ProductNode_POSIT9258: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2201Output_11459,ProductNode_POSIT2521Output_3119,ProductNode_POSIT9258Output_11460);

ProductNode_POSIT9267: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2203Output_11470,ProductNode_POSIT2524Output_3123,ProductNode_POSIT9267Output_11471);

ProductNode_POSIT9275: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2205Output_11480,ProductNode_POSIT2532Output_3133,ProductNode_POSIT9275Output_11481);

SumNode_POSIT2206: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT9275Output_11481,ProductNode_POSIT9267Output_11471,SumNode_POSIT2206Output_11482);

ProductNode_POSIT9276: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2206Output_11482,ProductNode_POSIT2539Output_3142,ProductNode_POSIT9276Output_11483);

SumNode_POSIT2207: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT9276Output_11483,ProductNode_POSIT9258Output_11460,SumNode_POSIT2207Output_11484);

ProductNode_POSIT9277: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2207Output_11484,ProductNode_POSIT9240Output_11437,ProductNode_POSIT9277Output_11485);

ProductNode_POSIT9304: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT9304weight,ProductNode_POSIT2583Output_3196,ProductNode_POSIT9304Output_11516);

ProductNode_POSIT9308: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT9308weight,ProductNode_POSIT2587Output_3201,ProductNode_POSIT9308Output_11521);

SumNode_POSIT2213: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT9308Output_11521,ProductNode_POSIT9304Output_11516,SumNode_POSIT2213Output_11522);

ProductNode_POSIT9309: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2213Output_11522,ProductNode_POSIT7621Output_9433,ProductNode_POSIT9309Output_11523);

ProductNode_POSIT9336: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT9336weight,ProductNode_POSIT2583Output_3196,ProductNode_POSIT9336Output_11554);

ProductNode_POSIT9340: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT9340weight,ProductNode_POSIT2587Output_3201,ProductNode_POSIT9340Output_11559);

SumNode_POSIT2219: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT9340Output_11559,ProductNode_POSIT9336Output_11554,SumNode_POSIT2219Output_11560);

ProductNode_POSIT9341: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2219Output_11560,ProductNode_POSIT7653Output_9471,ProductNode_POSIT9341Output_11561);

SumNode_POSIT2220: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT9341Output_11561,ProductNode_POSIT9309Output_11523,SumNode_POSIT2220Output_11562);

ProductNode_POSIT9342: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2220Output_11562,ProductNode_POSIT9277Output_11485,ProductNode_POSIT9342Output_11563);

ProductNode_POSIT9344: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT9344weight,ProductNode_POSIT2623Output_3245,ProductNode_POSIT9344Output_11565);

ProductNode_POSIT9353: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2222Output_11575,ProductNode_POSIT2524Output_3123,ProductNode_POSIT9353Output_11576);

ProductNode_POSIT9361: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2224Output_11585,ProductNode_POSIT2532Output_3133,ProductNode_POSIT9361Output_11586);

SumNode_POSIT2225: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT9361Output_11586,ProductNode_POSIT9353Output_11576,SumNode_POSIT2225Output_11587);

ProductNode_POSIT9362: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2225Output_11587,ProductNode_POSIT2521Output_3119,ProductNode_POSIT9362Output_11588);

ProductNode_POSIT9371: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2227Output_11598,ProductNode_POSIT2524Output_3123,ProductNode_POSIT9371Output_11599);

ProductNode_POSIT9379: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2229Output_11608,ProductNode_POSIT2532Output_3133,ProductNode_POSIT9379Output_11609);

SumNode_POSIT2230: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT9379Output_11609,ProductNode_POSIT9371Output_11599,SumNode_POSIT2230Output_11610);

ProductNode_POSIT9380: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2230Output_11610,ProductNode_POSIT2539Output_3142,ProductNode_POSIT9380Output_11611);

SumNode_POSIT2231: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT9380Output_11611,ProductNode_POSIT9362Output_11588,SumNode_POSIT2231Output_11612);

ProductNode_POSIT9381: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2231Output_11612,ProductNode_POSIT9344Output_11565,ProductNode_POSIT9381Output_11613);

ProductNode_POSIT9408: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT9408weight,ProductNode_POSIT2583Output_3196,ProductNode_POSIT9408Output_11644);

ProductNode_POSIT9412: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT9412weight,ProductNode_POSIT2587Output_3201,ProductNode_POSIT9412Output_11649);

SumNode_POSIT2237: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT9412Output_11649,ProductNode_POSIT9408Output_11644,SumNode_POSIT2237Output_11650);

ProductNode_POSIT9413: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2237Output_11650,ProductNode_POSIT7725Output_9561,ProductNode_POSIT9413Output_11651);

ProductNode_POSIT9440: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT9440weight,ProductNode_POSIT2583Output_3196,ProductNode_POSIT9440Output_11682);

ProductNode_POSIT9444: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT9444weight,ProductNode_POSIT2587Output_3201,ProductNode_POSIT9444Output_11687);

SumNode_POSIT2243: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT9444Output_11687,ProductNode_POSIT9440Output_11682,SumNode_POSIT2243Output_11688);

ProductNode_POSIT9445: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2243Output_11688,ProductNode_POSIT7757Output_9599,ProductNode_POSIT9445Output_11689);

SumNode_POSIT2244: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT9445Output_11689,ProductNode_POSIT9413Output_11651,SumNode_POSIT2244Output_11690);

ProductNode_POSIT9446: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2244Output_11690,ProductNode_POSIT9381Output_11613,ProductNode_POSIT9446Output_11691);

SumNode_POSIT2245: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT9446Output_11691,ProductNode_POSIT9342Output_11563,SumNode_POSIT2245Output_11692);

ProductNode_POSIT9447: entity work.PositMult_23_6_comb_uid2(arch)
port map(v13,SumNode_POSIT2245Output_11692,ProductNode_POSIT9447Output_11693);

ProductNode_POSIT9449: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT9449weight,ProductNode_POSIT2519Output_3117,ProductNode_POSIT9449Output_11695);

ProductNode_POSIT9486: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2256Output_11742,ProductNode_POSIT9449Output_11695,ProductNode_POSIT9486Output_11743);

ProductNode_POSIT9513: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT9513weight,ProductNode_POSIT2792Output_3454,ProductNode_POSIT9513Output_11774);

ProductNode_POSIT9517: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT9517weight,ProductNode_POSIT2796Output_3459,ProductNode_POSIT9517Output_11779);

SumNode_POSIT2262: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT9517Output_11779,ProductNode_POSIT9513Output_11774,SumNode_POSIT2262Output_11780);

ProductNode_POSIT9518: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2262Output_11780,ProductNode_POSIT7621Output_9433,ProductNode_POSIT9518Output_11781);

ProductNode_POSIT9545: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT9545weight,ProductNode_POSIT2792Output_3454,ProductNode_POSIT9545Output_11812);

ProductNode_POSIT9549: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT9549weight,ProductNode_POSIT2796Output_3459,ProductNode_POSIT9549Output_11817);

SumNode_POSIT2268: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT9549Output_11817,ProductNode_POSIT9545Output_11812,SumNode_POSIT2268Output_11818);

ProductNode_POSIT9550: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2268Output_11818,ProductNode_POSIT7653Output_9471,ProductNode_POSIT9550Output_11819);

SumNode_POSIT2269: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT9550Output_11819,ProductNode_POSIT9518Output_11781,SumNode_POSIT2269Output_11820);

ProductNode_POSIT9551: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2269Output_11820,ProductNode_POSIT9486Output_11743,ProductNode_POSIT9551Output_11821);

ProductNode_POSIT9553: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT9553weight,ProductNode_POSIT2623Output_3245,ProductNode_POSIT9553Output_11823);

ProductNode_POSIT9590: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2280Output_11870,ProductNode_POSIT9553Output_11823,ProductNode_POSIT9590Output_11871);

ProductNode_POSIT9617: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT9617weight,ProductNode_POSIT2792Output_3454,ProductNode_POSIT9617Output_11902);

ProductNode_POSIT9621: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT9621weight,ProductNode_POSIT2796Output_3459,ProductNode_POSIT9621Output_11907);

SumNode_POSIT2286: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT9621Output_11907,ProductNode_POSIT9617Output_11902,SumNode_POSIT2286Output_11908);

ProductNode_POSIT9622: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2286Output_11908,ProductNode_POSIT7725Output_9561,ProductNode_POSIT9622Output_11909);

ProductNode_POSIT9649: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT9649weight,ProductNode_POSIT2792Output_3454,ProductNode_POSIT9649Output_11940);

ProductNode_POSIT9653: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT9653weight,ProductNode_POSIT2796Output_3459,ProductNode_POSIT9653Output_11945);

SumNode_POSIT2292: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT9653Output_11945,ProductNode_POSIT9649Output_11940,SumNode_POSIT2292Output_11946);

ProductNode_POSIT9654: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2292Output_11946,ProductNode_POSIT7757Output_9599,ProductNode_POSIT9654Output_11947);

SumNode_POSIT2293: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT9654Output_11947,ProductNode_POSIT9622Output_11909,SumNode_POSIT2293Output_11948);

ProductNode_POSIT9655: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2293Output_11948,ProductNode_POSIT9590Output_11871,ProductNode_POSIT9655Output_11949);

SumNode_POSIT2294: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT9655Output_11949,ProductNode_POSIT9551Output_11821,SumNode_POSIT2294Output_11950);

ProductNode_POSIT9656: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb13,SumNode_POSIT2294Output_11950,ProductNode_POSIT9656Output_11951);

SumNode_POSIT2295: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT9656Output_11951,ProductNode_POSIT9447Output_11693,SumNode_POSIT2295Output_11952);

ProductNode_POSIT9657: entity work.PositMult_23_6_comb_uid2(arch)
port map(v3,SumNode_POSIT2295Output_11952,ProductNode_POSIT9657Output_11953);

ProductNode_POSIT9677: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2300Output_11977,ProductNode_POSIT2940Output_3637,ProductNode_POSIT9677Output_11978);

ProductNode_POSIT9695: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2305Output_12000,ProductNode_POSIT2958Output_3660,ProductNode_POSIT9695Output_12001);

SumNode_POSIT2306: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT9695Output_12001,ProductNode_POSIT9677Output_11978,SumNode_POSIT2306Output_12002);

ProductNode_POSIT9696: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2306Output_12002,ProductNode_POSIT9240Output_11437,ProductNode_POSIT9696Output_12003);

ProductNode_POSIT9723: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT9723weight,ProductNode_POSIT2583Output_3196,ProductNode_POSIT9723Output_12034);

ProductNode_POSIT9727: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT9727weight,ProductNode_POSIT2587Output_3201,ProductNode_POSIT9727Output_12039);

SumNode_POSIT2312: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT9727Output_12039,ProductNode_POSIT9723Output_12034,SumNode_POSIT2312Output_12040);

ProductNode_POSIT9728: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2312Output_12040,ProductNode_POSIT8040Output_9951,ProductNode_POSIT9728Output_12041);

ProductNode_POSIT9755: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT9755weight,ProductNode_POSIT2583Output_3196,ProductNode_POSIT9755Output_12072);

ProductNode_POSIT9759: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT9759weight,ProductNode_POSIT2587Output_3201,ProductNode_POSIT9759Output_12077);

SumNode_POSIT2318: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT9759Output_12077,ProductNode_POSIT9755Output_12072,SumNode_POSIT2318Output_12078);

ProductNode_POSIT9760: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2318Output_12078,ProductNode_POSIT8072Output_9989,ProductNode_POSIT9760Output_12079);

SumNode_POSIT2319: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT9760Output_12079,ProductNode_POSIT9728Output_12041,SumNode_POSIT2319Output_12080);

ProductNode_POSIT9761: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2319Output_12080,ProductNode_POSIT9696Output_12003,ProductNode_POSIT9761Output_12081);

ProductNode_POSIT9781: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2324Output_12105,ProductNode_POSIT2940Output_3637,ProductNode_POSIT9781Output_12106);

ProductNode_POSIT9799: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2329Output_12128,ProductNode_POSIT2958Output_3660,ProductNode_POSIT9799Output_12129);

SumNode_POSIT2330: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT9799Output_12129,ProductNode_POSIT9781Output_12106,SumNode_POSIT2330Output_12130);

ProductNode_POSIT9800: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2330Output_12130,ProductNode_POSIT9344Output_11565,ProductNode_POSIT9800Output_12131);

ProductNode_POSIT9827: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT9827weight,ProductNode_POSIT2583Output_3196,ProductNode_POSIT9827Output_12162);

ProductNode_POSIT9831: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT9831weight,ProductNode_POSIT2587Output_3201,ProductNode_POSIT9831Output_12167);

SumNode_POSIT2336: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT9831Output_12167,ProductNode_POSIT9827Output_12162,SumNode_POSIT2336Output_12168);

ProductNode_POSIT9832: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2336Output_12168,ProductNode_POSIT8144Output_10079,ProductNode_POSIT9832Output_12169);

ProductNode_POSIT9859: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT9859weight,ProductNode_POSIT2583Output_3196,ProductNode_POSIT9859Output_12200);

ProductNode_POSIT9863: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT9863weight,ProductNode_POSIT2587Output_3201,ProductNode_POSIT9863Output_12205);

SumNode_POSIT2342: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT9863Output_12205,ProductNode_POSIT9859Output_12200,SumNode_POSIT2342Output_12206);

ProductNode_POSIT9864: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2342Output_12206,ProductNode_POSIT8176Output_10117,ProductNode_POSIT9864Output_12207);

SumNode_POSIT2343: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT9864Output_12207,ProductNode_POSIT9832Output_12169,SumNode_POSIT2343Output_12208);

ProductNode_POSIT9865: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2343Output_12208,ProductNode_POSIT9800Output_12131,ProductNode_POSIT9865Output_12209);

SumNode_POSIT2344: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT9865Output_12209,ProductNode_POSIT9761Output_12081,SumNode_POSIT2344Output_12210);

ProductNode_POSIT9866: entity work.PositMult_23_6_comb_uid2(arch)
port map(v13,SumNode_POSIT2344Output_12210,ProductNode_POSIT9866Output_12211);

ProductNode_POSIT9905: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2355Output_12260,ProductNode_POSIT9449Output_11695,ProductNode_POSIT9905Output_12261);

ProductNode_POSIT9932: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT9932weight,ProductNode_POSIT2792Output_3454,ProductNode_POSIT9932Output_12292);

ProductNode_POSIT9936: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT9936weight,ProductNode_POSIT2796Output_3459,ProductNode_POSIT9936Output_12297);

SumNode_POSIT2361: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT9936Output_12297,ProductNode_POSIT9932Output_12292,SumNode_POSIT2361Output_12298);

ProductNode_POSIT9937: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2361Output_12298,ProductNode_POSIT8040Output_9951,ProductNode_POSIT9937Output_12299);

ProductNode_POSIT9964: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT9964weight,ProductNode_POSIT2792Output_3454,ProductNode_POSIT9964Output_12330);

ProductNode_POSIT9968: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT9968weight,ProductNode_POSIT2796Output_3459,ProductNode_POSIT9968Output_12335);

SumNode_POSIT2367: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT9968Output_12335,ProductNode_POSIT9964Output_12330,SumNode_POSIT2367Output_12336);

ProductNode_POSIT9969: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2367Output_12336,ProductNode_POSIT8072Output_9989,ProductNode_POSIT9969Output_12337);

SumNode_POSIT2368: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT9969Output_12337,ProductNode_POSIT9937Output_12299,SumNode_POSIT2368Output_12338);

ProductNode_POSIT9970: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2368Output_12338,ProductNode_POSIT9905Output_12261,ProductNode_POSIT9970Output_12339);

ProductNode_POSIT10009: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2379Output_12388,ProductNode_POSIT9553Output_11823,ProductNode_POSIT10009Output_12389);

ProductNode_POSIT10036: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT10036weight,ProductNode_POSIT2792Output_3454,ProductNode_POSIT10036Output_12420);

ProductNode_POSIT10040: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT10040weight,ProductNode_POSIT2796Output_3459,ProductNode_POSIT10040Output_12425);

SumNode_POSIT2385: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT10040Output_12425,ProductNode_POSIT10036Output_12420,SumNode_POSIT2385Output_12426);

ProductNode_POSIT10041: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2385Output_12426,ProductNode_POSIT8144Output_10079,ProductNode_POSIT10041Output_12427);

ProductNode_POSIT10068: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT10068weight,ProductNode_POSIT2792Output_3454,ProductNode_POSIT10068Output_12458);

ProductNode_POSIT10072: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT10072weight,ProductNode_POSIT2796Output_3459,ProductNode_POSIT10072Output_12463);

SumNode_POSIT2391: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT10072Output_12463,ProductNode_POSIT10068Output_12458,SumNode_POSIT2391Output_12464);

ProductNode_POSIT10073: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2391Output_12464,ProductNode_POSIT8176Output_10117,ProductNode_POSIT10073Output_12465);

SumNode_POSIT2392: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT10073Output_12465,ProductNode_POSIT10041Output_12427,SumNode_POSIT2392Output_12466);

ProductNode_POSIT10074: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2392Output_12466,ProductNode_POSIT10009Output_12389,ProductNode_POSIT10074Output_12467);

SumNode_POSIT2393: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT10074Output_12467,ProductNode_POSIT9970Output_12339,SumNode_POSIT2393Output_12468);

ProductNode_POSIT10075: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb13,SumNode_POSIT2393Output_12468,ProductNode_POSIT10075Output_12469);

SumNode_POSIT2394: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT10075Output_12469,ProductNode_POSIT9866Output_12211,SumNode_POSIT2394Output_12470);

ProductNode_POSIT10076: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb3,SumNode_POSIT2394Output_12470,ProductNode_POSIT10076Output_12471);

SumNode_POSIT2395: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT10076Output_12471,ProductNode_POSIT9657Output_11953,SumNode_POSIT2395Output_12472);

ProductNode_POSIT10077: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb4,SumNode_POSIT2395Output_12472,ProductNode_POSIT10077Output_12473);

SumNode_POSIT2396: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT10077Output_12473,ProductNode_POSIT9238Output_11435,SumNode_POSIT2396Output_12474);

ProductNode_POSIT10078: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb12,SumNode_POSIT2396Output_12474,ProductNode_POSIT10078Output_12475);

SumNode_POSIT2397: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT10078Output_12475,ProductNode_POSIT8399Output_10397,SumNode_POSIT2397Output_12476);

ProductNode_POSIT10079: entity work.PositMult_23_6_comb_uid2(arch)
port map(v6,SumNode_POSIT2397Output_12476,ProductNode_POSIT10079Output_12477);

ProductNode_POSIT10081: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT10081weight,ProductNode_POSIT1Output_1,ProductNode_POSIT10081Output_12479);

ProductNode_POSIT10090: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2399Output_12489,ProductNode_POSIT3365Output_4165,ProductNode_POSIT10090Output_12490);

ProductNode_POSIT10098: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2401Output_12499,ProductNode_POSIT3373Output_4175,ProductNode_POSIT10098Output_12500);

SumNode_POSIT2402: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT10098Output_12500,ProductNode_POSIT10090Output_12490,SumNode_POSIT2402Output_12501);

ProductNode_POSIT10099: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2402Output_12501,ProductNode_POSIT3Output_3,ProductNode_POSIT10099Output_12502);

ProductNode_POSIT10108: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2404Output_12512,ProductNode_POSIT3365Output_4165,ProductNode_POSIT10108Output_12513);

ProductNode_POSIT10116: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2406Output_12522,ProductNode_POSIT3373Output_4175,ProductNode_POSIT10116Output_12523);

SumNode_POSIT2407: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT10116Output_12523,ProductNode_POSIT10108Output_12513,SumNode_POSIT2407Output_12524);

ProductNode_POSIT10117: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2407Output_12524,ProductNode_POSIT21Output_26,ProductNode_POSIT10117Output_12525);

SumNode_POSIT2408: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT10117Output_12525,ProductNode_POSIT10099Output_12502,SumNode_POSIT2408Output_12526);

ProductNode_POSIT10118: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2408Output_12526,ProductNode_POSIT10081Output_12479,ProductNode_POSIT10118Output_12527);

ProductNode_POSIT10140: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT812Output_4232,ProductNode_POSIT6760Output_8370,ProductNode_POSIT10140Output_12552);

ProductNode_POSIT10141: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT10141weight,ProductNode_POSIT10140Output_12552,ProductNode_POSIT10141Output_12553);

ProductNode_POSIT10150: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2414Output_12564,ProductNode_POSIT10141Output_12553,ProductNode_POSIT10150Output_12565);

ProductNode_POSIT10172: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT818Output_4270,ProductNode_POSIT6792Output_8408,ProductNode_POSIT10172Output_12590);

ProductNode_POSIT10173: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT10173weight,ProductNode_POSIT10172Output_12590,ProductNode_POSIT10173Output_12591);

ProductNode_POSIT10182: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2420Output_12602,ProductNode_POSIT10173Output_12591,ProductNode_POSIT10182Output_12603);

SumNode_POSIT2421: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT10182Output_12603,ProductNode_POSIT10150Output_12565,SumNode_POSIT2421Output_12604);

ProductNode_POSIT10183: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2421Output_12604,ProductNode_POSIT10118Output_12527,ProductNode_POSIT10183Output_12605);

ProductNode_POSIT10185: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT10185weight,ProductNode_POSIT105Output_129,ProductNode_POSIT10185Output_12607);

ProductNode_POSIT10194: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2423Output_12617,ProductNode_POSIT3365Output_4165,ProductNode_POSIT10194Output_12618);

ProductNode_POSIT10202: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2425Output_12627,ProductNode_POSIT3373Output_4175,ProductNode_POSIT10202Output_12628);

SumNode_POSIT2426: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT10202Output_12628,ProductNode_POSIT10194Output_12618,SumNode_POSIT2426Output_12629);

ProductNode_POSIT10203: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2426Output_12629,ProductNode_POSIT3Output_3,ProductNode_POSIT10203Output_12630);

ProductNode_POSIT10212: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2428Output_12640,ProductNode_POSIT3365Output_4165,ProductNode_POSIT10212Output_12641);

ProductNode_POSIT10220: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2430Output_12650,ProductNode_POSIT3373Output_4175,ProductNode_POSIT10220Output_12651);

SumNode_POSIT2431: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT10220Output_12651,ProductNode_POSIT10212Output_12641,SumNode_POSIT2431Output_12652);

ProductNode_POSIT10221: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2431Output_12652,ProductNode_POSIT21Output_26,ProductNode_POSIT10221Output_12653);

SumNode_POSIT2432: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT10221Output_12653,ProductNode_POSIT10203Output_12630,SumNode_POSIT2432Output_12654);

ProductNode_POSIT10222: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2432Output_12654,ProductNode_POSIT10185Output_12607,ProductNode_POSIT10222Output_12655);

ProductNode_POSIT10245: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT10245weight,ProductNode_POSIT10140Output_12552,ProductNode_POSIT10245Output_12681);

ProductNode_POSIT10254: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2438Output_12692,ProductNode_POSIT10245Output_12681,ProductNode_POSIT10254Output_12693);

ProductNode_POSIT10277: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT10277weight,ProductNode_POSIT10172Output_12590,ProductNode_POSIT10277Output_12719);

ProductNode_POSIT10286: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2444Output_12730,ProductNode_POSIT10277Output_12719,ProductNode_POSIT10286Output_12731);

SumNode_POSIT2445: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT10286Output_12731,ProductNode_POSIT10254Output_12693,SumNode_POSIT2445Output_12732);

ProductNode_POSIT10287: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2445Output_12732,ProductNode_POSIT10222Output_12655,ProductNode_POSIT10287Output_12733);

SumNode_POSIT2446: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT10287Output_12733,ProductNode_POSIT10183Output_12605,SumNode_POSIT2446Output_12734);

ProductNode_POSIT10288: entity work.PositMult_23_6_comb_uid2(arch)
port map(v13,SumNode_POSIT2446Output_12734,ProductNode_POSIT10288Output_12735);

ProductNode_POSIT10290: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT10290weight,ProductNode_POSIT1Output_1,ProductNode_POSIT10290Output_12737);

ProductNode_POSIT10327: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2457Output_12784,ProductNode_POSIT10290Output_12737,ProductNode_POSIT10327Output_12785);

ProductNode_POSIT10359: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1664Output_8664,ProductNode_POSIT10141Output_12553,ProductNode_POSIT10359Output_12823);

ProductNode_POSIT10391: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1670Output_8702,ProductNode_POSIT10173Output_12591,ProductNode_POSIT10391Output_12861);

SumNode_POSIT2470: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT10391Output_12861,ProductNode_POSIT10359Output_12823,SumNode_POSIT2470Output_12862);

ProductNode_POSIT10392: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2470Output_12862,ProductNode_POSIT10327Output_12785,ProductNode_POSIT10392Output_12863);

ProductNode_POSIT10394: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT10394weight,ProductNode_POSIT105Output_129,ProductNode_POSIT10394Output_12865);

ProductNode_POSIT10431: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2481Output_12912,ProductNode_POSIT10394Output_12865,ProductNode_POSIT10431Output_12913);

ProductNode_POSIT10463: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1688Output_8792,ProductNode_POSIT10245Output_12681,ProductNode_POSIT10463Output_12951);

ProductNode_POSIT10495: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1694Output_8830,ProductNode_POSIT10277Output_12719,ProductNode_POSIT10495Output_12989);

SumNode_POSIT2494: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT10495Output_12989,ProductNode_POSIT10463Output_12951,SumNode_POSIT2494Output_12990);

ProductNode_POSIT10496: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2494Output_12990,ProductNode_POSIT10431Output_12913,ProductNode_POSIT10496Output_12991);

SumNode_POSIT2495: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT10496Output_12991,ProductNode_POSIT10392Output_12863,SumNode_POSIT2495Output_12992);

ProductNode_POSIT10497: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb13,SumNode_POSIT2495Output_12992,ProductNode_POSIT10497Output_12993);

SumNode_POSIT2496: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT10497Output_12993,ProductNode_POSIT10288Output_12735,SumNode_POSIT2496Output_12994);

ProductNode_POSIT10498: entity work.PositMult_23_6_comb_uid2(arch)
port map(v3,SumNode_POSIT2496Output_12994,ProductNode_POSIT10498Output_12995);

ProductNode_POSIT10518: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2501Output_13019,ProductNode_POSIT422Output_521,ProductNode_POSIT10518Output_13020);

ProductNode_POSIT10536: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2506Output_13042,ProductNode_POSIT440Output_544,ProductNode_POSIT10536Output_13043);

SumNode_POSIT2507: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT10536Output_13043,ProductNode_POSIT10518Output_13020,SumNode_POSIT2507Output_13044);

ProductNode_POSIT10537: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2507Output_13044,ProductNode_POSIT10081Output_12479,ProductNode_POSIT10537Output_13045);

ProductNode_POSIT10559: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT911Output_4750,ProductNode_POSIT6760Output_8370,ProductNode_POSIT10559Output_13070);

ProductNode_POSIT10560: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT10560weight,ProductNode_POSIT10559Output_13070,ProductNode_POSIT10560Output_13071);

ProductNode_POSIT10569: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2513Output_13082,ProductNode_POSIT10560Output_13071,ProductNode_POSIT10569Output_13083);

ProductNode_POSIT10591: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT917Output_4788,ProductNode_POSIT6792Output_8408,ProductNode_POSIT10591Output_13108);

ProductNode_POSIT10592: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT10592weight,ProductNode_POSIT10591Output_13108,ProductNode_POSIT10592Output_13109);

ProductNode_POSIT10601: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2519Output_13120,ProductNode_POSIT10592Output_13109,ProductNode_POSIT10601Output_13121);

SumNode_POSIT2520: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT10601Output_13121,ProductNode_POSIT10569Output_13083,SumNode_POSIT2520Output_13122);

ProductNode_POSIT10602: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2520Output_13122,ProductNode_POSIT10537Output_13045,ProductNode_POSIT10602Output_13123);

ProductNode_POSIT10622: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2525Output_13147,ProductNode_POSIT422Output_521,ProductNode_POSIT10622Output_13148);

ProductNode_POSIT10640: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2530Output_13170,ProductNode_POSIT440Output_544,ProductNode_POSIT10640Output_13171);

SumNode_POSIT2531: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT10640Output_13171,ProductNode_POSIT10622Output_13148,SumNode_POSIT2531Output_13172);

ProductNode_POSIT10641: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2531Output_13172,ProductNode_POSIT10185Output_12607,ProductNode_POSIT10641Output_13173);

ProductNode_POSIT10664: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT10664weight,ProductNode_POSIT10559Output_13070,ProductNode_POSIT10664Output_13199);

ProductNode_POSIT10673: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2537Output_13210,ProductNode_POSIT10664Output_13199,ProductNode_POSIT10673Output_13211);

ProductNode_POSIT10696: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT10696weight,ProductNode_POSIT10591Output_13108,ProductNode_POSIT10696Output_13237);

ProductNode_POSIT10705: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2543Output_13248,ProductNode_POSIT10696Output_13237,ProductNode_POSIT10705Output_13249);

SumNode_POSIT2544: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT10705Output_13249,ProductNode_POSIT10673Output_13211,SumNode_POSIT2544Output_13250);

ProductNode_POSIT10706: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2544Output_13250,ProductNode_POSIT10641Output_13173,ProductNode_POSIT10706Output_13251);

SumNode_POSIT2545: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT10706Output_13251,ProductNode_POSIT10602Output_13123,SumNode_POSIT2545Output_13252);

ProductNode_POSIT10707: entity work.PositMult_23_6_comb_uid2(arch)
port map(v13,SumNode_POSIT2545Output_13252,ProductNode_POSIT10707Output_13253);

ProductNode_POSIT10746: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2556Output_13302,ProductNode_POSIT10290Output_12737,ProductNode_POSIT10746Output_13303);

ProductNode_POSIT10778: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1763Output_9182,ProductNode_POSIT10560Output_13071,ProductNode_POSIT10778Output_13341);

ProductNode_POSIT10810: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1769Output_9220,ProductNode_POSIT10592Output_13109,ProductNode_POSIT10810Output_13379);

SumNode_POSIT2569: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT10810Output_13379,ProductNode_POSIT10778Output_13341,SumNode_POSIT2569Output_13380);

ProductNode_POSIT10811: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2569Output_13380,ProductNode_POSIT10746Output_13303,ProductNode_POSIT10811Output_13381);

ProductNode_POSIT10850: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2580Output_13430,ProductNode_POSIT10394Output_12865,ProductNode_POSIT10850Output_13431);

ProductNode_POSIT10882: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1787Output_9310,ProductNode_POSIT10664Output_13199,ProductNode_POSIT10882Output_13469);

ProductNode_POSIT10914: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1793Output_9348,ProductNode_POSIT10696Output_13237,ProductNode_POSIT10914Output_13507);

SumNode_POSIT2593: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT10914Output_13507,ProductNode_POSIT10882Output_13469,SumNode_POSIT2593Output_13508);

ProductNode_POSIT10915: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2593Output_13508,ProductNode_POSIT10850Output_13431,ProductNode_POSIT10915Output_13509);

SumNode_POSIT2594: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT10915Output_13509,ProductNode_POSIT10811Output_13381,SumNode_POSIT2594Output_13510);

ProductNode_POSIT10916: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb13,SumNode_POSIT2594Output_13510,ProductNode_POSIT10916Output_13511);

SumNode_POSIT2595: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT10916Output_13511,ProductNode_POSIT10707Output_13253,SumNode_POSIT2595Output_13512);

ProductNode_POSIT10917: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb3,SumNode_POSIT2595Output_13512,ProductNode_POSIT10917Output_13513);

SumNode_POSIT2596: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT10917Output_13513,ProductNode_POSIT10498Output_12995,SumNode_POSIT2596Output_13514);

ProductNode_POSIT10918: entity work.PositMult_23_6_comb_uid2(arch)
port map(v4,SumNode_POSIT2596Output_13514,ProductNode_POSIT10918Output_13515);

ProductNode_POSIT10920: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT10920weight,ProductNode_POSIT840Output_1039,ProductNode_POSIT10920Output_13517);

ProductNode_POSIT10929: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2598Output_13527,ProductNode_POSIT4204Output_5203,ProductNode_POSIT10929Output_13528);

ProductNode_POSIT10937: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2600Output_13537,ProductNode_POSIT4212Output_5213,ProductNode_POSIT10937Output_13538);

SumNode_POSIT2601: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT10937Output_13538,ProductNode_POSIT10929Output_13528,SumNode_POSIT2601Output_13539);

ProductNode_POSIT10938: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2601Output_13539,ProductNode_POSIT842Output_1041,ProductNode_POSIT10938Output_13540);

ProductNode_POSIT10947: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2603Output_13550,ProductNode_POSIT4204Output_5203,ProductNode_POSIT10947Output_13551);

ProductNode_POSIT10955: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2605Output_13560,ProductNode_POSIT4212Output_5213,ProductNode_POSIT10955Output_13561);

SumNode_POSIT2606: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT10955Output_13561,ProductNode_POSIT10947Output_13551,SumNode_POSIT2606Output_13562);

ProductNode_POSIT10956: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2606Output_13562,ProductNode_POSIT860Output_1064,ProductNode_POSIT10956Output_13563);

SumNode_POSIT2607: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT10956Output_13563,ProductNode_POSIT10938Output_13540,SumNode_POSIT2607Output_13564);

ProductNode_POSIT10957: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2607Output_13564,ProductNode_POSIT10920Output_13517,ProductNode_POSIT10957Output_13565);

ProductNode_POSIT10979: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1011Output_5270,ProductNode_POSIT6760Output_8370,ProductNode_POSIT10979Output_13590);

ProductNode_POSIT10980: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT10980weight,ProductNode_POSIT10979Output_13590,ProductNode_POSIT10980Output_13591);

ProductNode_POSIT10989: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2613Output_13602,ProductNode_POSIT10980Output_13591,ProductNode_POSIT10989Output_13603);

ProductNode_POSIT11011: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1017Output_5308,ProductNode_POSIT6792Output_8408,ProductNode_POSIT11011Output_13628);

ProductNode_POSIT11012: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT11012weight,ProductNode_POSIT11011Output_13628,ProductNode_POSIT11012Output_13629);

ProductNode_POSIT11021: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2619Output_13640,ProductNode_POSIT11012Output_13629,ProductNode_POSIT11021Output_13641);

SumNode_POSIT2620: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT11021Output_13641,ProductNode_POSIT10989Output_13603,SumNode_POSIT2620Output_13642);

ProductNode_POSIT11022: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2620Output_13642,ProductNode_POSIT10957Output_13565,ProductNode_POSIT11022Output_13643);

ProductNode_POSIT11024: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT11024weight,ProductNode_POSIT944Output_1167,ProductNode_POSIT11024Output_13645);

ProductNode_POSIT11033: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2622Output_13655,ProductNode_POSIT4204Output_5203,ProductNode_POSIT11033Output_13656);

ProductNode_POSIT11041: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2624Output_13665,ProductNode_POSIT4212Output_5213,ProductNode_POSIT11041Output_13666);

SumNode_POSIT2625: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT11041Output_13666,ProductNode_POSIT11033Output_13656,SumNode_POSIT2625Output_13667);

ProductNode_POSIT11042: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2625Output_13667,ProductNode_POSIT842Output_1041,ProductNode_POSIT11042Output_13668);

ProductNode_POSIT11051: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2627Output_13678,ProductNode_POSIT4204Output_5203,ProductNode_POSIT11051Output_13679);

ProductNode_POSIT11059: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2629Output_13688,ProductNode_POSIT4212Output_5213,ProductNode_POSIT11059Output_13689);

SumNode_POSIT2630: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT11059Output_13689,ProductNode_POSIT11051Output_13679,SumNode_POSIT2630Output_13690);

ProductNode_POSIT11060: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2630Output_13690,ProductNode_POSIT860Output_1064,ProductNode_POSIT11060Output_13691);

SumNode_POSIT2631: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT11060Output_13691,ProductNode_POSIT11042Output_13668,SumNode_POSIT2631Output_13692);

ProductNode_POSIT11061: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2631Output_13692,ProductNode_POSIT11024Output_13645,ProductNode_POSIT11061Output_13693);

ProductNode_POSIT11084: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT11084weight,ProductNode_POSIT10979Output_13590,ProductNode_POSIT11084Output_13719);

ProductNode_POSIT11093: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2637Output_13730,ProductNode_POSIT11084Output_13719,ProductNode_POSIT11093Output_13731);

ProductNode_POSIT11116: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT11116weight,ProductNode_POSIT11011Output_13628,ProductNode_POSIT11116Output_13757);

ProductNode_POSIT11125: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2643Output_13768,ProductNode_POSIT11116Output_13757,ProductNode_POSIT11125Output_13769);

SumNode_POSIT2644: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT11125Output_13769,ProductNode_POSIT11093Output_13731,SumNode_POSIT2644Output_13770);

ProductNode_POSIT11126: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2644Output_13770,ProductNode_POSIT11061Output_13693,ProductNode_POSIT11126Output_13771);

SumNode_POSIT2645: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT11126Output_13771,ProductNode_POSIT11022Output_13643,SumNode_POSIT2645Output_13772);

ProductNode_POSIT11127: entity work.PositMult_23_6_comb_uid2(arch)
port map(v13,SumNode_POSIT2645Output_13772,ProductNode_POSIT11127Output_13773);

ProductNode_POSIT11129: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT11129weight,ProductNode_POSIT840Output_1039,ProductNode_POSIT11129Output_13775);

ProductNode_POSIT11166: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2656Output_13822,ProductNode_POSIT11129Output_13775,ProductNode_POSIT11166Output_13823);

ProductNode_POSIT11198: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1863Output_9702,ProductNode_POSIT10980Output_13591,ProductNode_POSIT11198Output_13861);

ProductNode_POSIT11230: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1869Output_9740,ProductNode_POSIT11012Output_13629,ProductNode_POSIT11230Output_13899);

SumNode_POSIT2669: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT11230Output_13899,ProductNode_POSIT11198Output_13861,SumNode_POSIT2669Output_13900);

ProductNode_POSIT11231: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2669Output_13900,ProductNode_POSIT11166Output_13823,ProductNode_POSIT11231Output_13901);

ProductNode_POSIT11233: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT11233weight,ProductNode_POSIT944Output_1167,ProductNode_POSIT11233Output_13903);

ProductNode_POSIT11270: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2680Output_13950,ProductNode_POSIT11233Output_13903,ProductNode_POSIT11270Output_13951);

ProductNode_POSIT11302: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1887Output_9830,ProductNode_POSIT11084Output_13719,ProductNode_POSIT11302Output_13989);

ProductNode_POSIT11334: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1893Output_9868,ProductNode_POSIT11116Output_13757,ProductNode_POSIT11334Output_14027);

SumNode_POSIT2693: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT11334Output_14027,ProductNode_POSIT11302Output_13989,SumNode_POSIT2693Output_14028);

ProductNode_POSIT11335: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2693Output_14028,ProductNode_POSIT11270Output_13951,ProductNode_POSIT11335Output_14029);

SumNode_POSIT2694: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT11335Output_14029,ProductNode_POSIT11231Output_13901,SumNode_POSIT2694Output_14030);

ProductNode_POSIT11336: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb13,SumNode_POSIT2694Output_14030,ProductNode_POSIT11336Output_14031);

SumNode_POSIT2695: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT11336Output_14031,ProductNode_POSIT11127Output_13773,SumNode_POSIT2695Output_14032);

ProductNode_POSIT11337: entity work.PositMult_23_6_comb_uid2(arch)
port map(v3,SumNode_POSIT2695Output_14032,ProductNode_POSIT11337Output_14033);

ProductNode_POSIT11357: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2700Output_14057,ProductNode_POSIT1261Output_1559,ProductNode_POSIT11357Output_14058);

ProductNode_POSIT11375: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2705Output_14080,ProductNode_POSIT1279Output_1582,ProductNode_POSIT11375Output_14081);

SumNode_POSIT2706: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT11375Output_14081,ProductNode_POSIT11357Output_14058,SumNode_POSIT2706Output_14082);

ProductNode_POSIT11376: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2706Output_14082,ProductNode_POSIT10920Output_13517,ProductNode_POSIT11376Output_14083);

ProductNode_POSIT11398: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1110Output_5788,ProductNode_POSIT6760Output_8370,ProductNode_POSIT11398Output_14108);

ProductNode_POSIT11399: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT11399weight,ProductNode_POSIT11398Output_14108,ProductNode_POSIT11399Output_14109);

ProductNode_POSIT11408: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2712Output_14120,ProductNode_POSIT11399Output_14109,ProductNode_POSIT11408Output_14121);

ProductNode_POSIT11430: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1116Output_5826,ProductNode_POSIT6792Output_8408,ProductNode_POSIT11430Output_14146);

ProductNode_POSIT11431: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT11431weight,ProductNode_POSIT11430Output_14146,ProductNode_POSIT11431Output_14147);

ProductNode_POSIT11440: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2718Output_14158,ProductNode_POSIT11431Output_14147,ProductNode_POSIT11440Output_14159);

SumNode_POSIT2719: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT11440Output_14159,ProductNode_POSIT11408Output_14121,SumNode_POSIT2719Output_14160);

ProductNode_POSIT11441: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2719Output_14160,ProductNode_POSIT11376Output_14083,ProductNode_POSIT11441Output_14161);

ProductNode_POSIT11461: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2724Output_14185,ProductNode_POSIT1261Output_1559,ProductNode_POSIT11461Output_14186);

ProductNode_POSIT11479: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2729Output_14208,ProductNode_POSIT1279Output_1582,ProductNode_POSIT11479Output_14209);

SumNode_POSIT2730: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT11479Output_14209,ProductNode_POSIT11461Output_14186,SumNode_POSIT2730Output_14210);

ProductNode_POSIT11480: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2730Output_14210,ProductNode_POSIT11024Output_13645,ProductNode_POSIT11480Output_14211);

ProductNode_POSIT11503: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT11503weight,ProductNode_POSIT11398Output_14108,ProductNode_POSIT11503Output_14237);

ProductNode_POSIT11512: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2736Output_14248,ProductNode_POSIT11503Output_14237,ProductNode_POSIT11512Output_14249);

ProductNode_POSIT11535: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT11535weight,ProductNode_POSIT11430Output_14146,ProductNode_POSIT11535Output_14275);

ProductNode_POSIT11544: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2742Output_14286,ProductNode_POSIT11535Output_14275,ProductNode_POSIT11544Output_14287);

SumNode_POSIT2743: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT11544Output_14287,ProductNode_POSIT11512Output_14249,SumNode_POSIT2743Output_14288);

ProductNode_POSIT11545: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2743Output_14288,ProductNode_POSIT11480Output_14211,ProductNode_POSIT11545Output_14289);

SumNode_POSIT2744: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT11545Output_14289,ProductNode_POSIT11441Output_14161,SumNode_POSIT2744Output_14290);

ProductNode_POSIT11546: entity work.PositMult_23_6_comb_uid2(arch)
port map(v13,SumNode_POSIT2744Output_14290,ProductNode_POSIT11546Output_14291);

ProductNode_POSIT11585: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2755Output_14340,ProductNode_POSIT11129Output_13775,ProductNode_POSIT11585Output_14341);

ProductNode_POSIT11617: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1962Output_10220,ProductNode_POSIT11399Output_14109,ProductNode_POSIT11617Output_14379);

ProductNode_POSIT11649: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1968Output_10258,ProductNode_POSIT11431Output_14147,ProductNode_POSIT11649Output_14417);

SumNode_POSIT2768: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT11649Output_14417,ProductNode_POSIT11617Output_14379,SumNode_POSIT2768Output_14418);

ProductNode_POSIT11650: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2768Output_14418,ProductNode_POSIT11585Output_14341,ProductNode_POSIT11650Output_14419);

ProductNode_POSIT11689: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2779Output_14468,ProductNode_POSIT11233Output_13903,ProductNode_POSIT11689Output_14469);

ProductNode_POSIT11721: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1986Output_10348,ProductNode_POSIT11503Output_14237,ProductNode_POSIT11721Output_14507);

ProductNode_POSIT11753: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT1992Output_10386,ProductNode_POSIT11535Output_14275,ProductNode_POSIT11753Output_14545);

SumNode_POSIT2792: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT11753Output_14545,ProductNode_POSIT11721Output_14507,SumNode_POSIT2792Output_14546);

ProductNode_POSIT11754: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2792Output_14546,ProductNode_POSIT11689Output_14469,ProductNode_POSIT11754Output_14547);

SumNode_POSIT2793: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT11754Output_14547,ProductNode_POSIT11650Output_14419,SumNode_POSIT2793Output_14548);

ProductNode_POSIT11755: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb13,SumNode_POSIT2793Output_14548,ProductNode_POSIT11755Output_14549);

SumNode_POSIT2794: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT11755Output_14549,ProductNode_POSIT11546Output_14291,SumNode_POSIT2794Output_14550);

ProductNode_POSIT11756: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb3,SumNode_POSIT2794Output_14550,ProductNode_POSIT11756Output_14551);

SumNode_POSIT2795: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT11756Output_14551,ProductNode_POSIT11337Output_14033,SumNode_POSIT2795Output_14552);

ProductNode_POSIT11757: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb4,SumNode_POSIT2795Output_14552,ProductNode_POSIT11757Output_14553);

SumNode_POSIT2796: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT11757Output_14553,ProductNode_POSIT10918Output_13515,SumNode_POSIT2796Output_14554);

ProductNode_POSIT11758: entity work.PositMult_23_6_comb_uid2(arch)
port map(v12,SumNode_POSIT2796Output_14554,ProductNode_POSIT11758Output_14555);

ProductNode_POSIT11760: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT11760weight,ProductNode_POSIT1680Output_2079,ProductNode_POSIT11760Output_14557);

ProductNode_POSIT11769: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2798Output_14567,ProductNode_POSIT5044Output_6243,ProductNode_POSIT11769Output_14568);

ProductNode_POSIT11777: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2800Output_14577,ProductNode_POSIT5052Output_6253,ProductNode_POSIT11777Output_14578);

SumNode_POSIT2801: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT11777Output_14578,ProductNode_POSIT11769Output_14568,SumNode_POSIT2801Output_14579);

ProductNode_POSIT11778: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2801Output_14579,ProductNode_POSIT1682Output_2081,ProductNode_POSIT11778Output_14580);

ProductNode_POSIT11787: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2803Output_14590,ProductNode_POSIT5044Output_6243,ProductNode_POSIT11787Output_14591);

ProductNode_POSIT11795: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2805Output_14600,ProductNode_POSIT5052Output_6253,ProductNode_POSIT11795Output_14601);

SumNode_POSIT2806: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT11795Output_14601,ProductNode_POSIT11787Output_14591,SumNode_POSIT2806Output_14602);

ProductNode_POSIT11796: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2806Output_14602,ProductNode_POSIT1700Output_2104,ProductNode_POSIT11796Output_14603);

SumNode_POSIT2807: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT11796Output_14603,ProductNode_POSIT11778Output_14580,SumNode_POSIT2807Output_14604);

ProductNode_POSIT11797: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2807Output_14604,ProductNode_POSIT11760Output_14557,ProductNode_POSIT11797Output_14605);

ProductNode_POSIT11829: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2014Output_10484,ProductNode_POSIT10141Output_12553,ProductNode_POSIT11829Output_14643);

ProductNode_POSIT11861: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2020Output_10522,ProductNode_POSIT10173Output_12591,ProductNode_POSIT11861Output_14681);

SumNode_POSIT2820: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT11861Output_14681,ProductNode_POSIT11829Output_14643,SumNode_POSIT2820Output_14682);

ProductNode_POSIT11862: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2820Output_14682,ProductNode_POSIT11797Output_14605,ProductNode_POSIT11862Output_14683);

ProductNode_POSIT11864: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT11864weight,ProductNode_POSIT1784Output_2207,ProductNode_POSIT11864Output_14685);

ProductNode_POSIT11873: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2822Output_14695,ProductNode_POSIT5044Output_6243,ProductNode_POSIT11873Output_14696);

ProductNode_POSIT11881: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2824Output_14705,ProductNode_POSIT5052Output_6253,ProductNode_POSIT11881Output_14706);

SumNode_POSIT2825: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT11881Output_14706,ProductNode_POSIT11873Output_14696,SumNode_POSIT2825Output_14707);

ProductNode_POSIT11882: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2825Output_14707,ProductNode_POSIT1682Output_2081,ProductNode_POSIT11882Output_14708);

ProductNode_POSIT11891: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2827Output_14718,ProductNode_POSIT5044Output_6243,ProductNode_POSIT11891Output_14719);

ProductNode_POSIT11899: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2829Output_14728,ProductNode_POSIT5052Output_6253,ProductNode_POSIT11899Output_14729);

SumNode_POSIT2830: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT11899Output_14729,ProductNode_POSIT11891Output_14719,SumNode_POSIT2830Output_14730);

ProductNode_POSIT11900: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2830Output_14730,ProductNode_POSIT1700Output_2104,ProductNode_POSIT11900Output_14731);

SumNode_POSIT2831: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT11900Output_14731,ProductNode_POSIT11882Output_14708,SumNode_POSIT2831Output_14732);

ProductNode_POSIT11901: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2831Output_14732,ProductNode_POSIT11864Output_14685,ProductNode_POSIT11901Output_14733);

ProductNode_POSIT11933: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2038Output_10612,ProductNode_POSIT10245Output_12681,ProductNode_POSIT11933Output_14771);

ProductNode_POSIT11965: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2044Output_10650,ProductNode_POSIT10277Output_12719,ProductNode_POSIT11965Output_14809);

SumNode_POSIT2844: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT11965Output_14809,ProductNode_POSIT11933Output_14771,SumNode_POSIT2844Output_14810);

ProductNode_POSIT11966: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2844Output_14810,ProductNode_POSIT11901Output_14733,ProductNode_POSIT11966Output_14811);

SumNode_POSIT2845: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT11966Output_14811,ProductNode_POSIT11862Output_14683,SumNode_POSIT2845Output_14812);

ProductNode_POSIT11967: entity work.PositMult_23_6_comb_uid2(arch)
port map(v13,SumNode_POSIT2845Output_14812,ProductNode_POSIT11967Output_14813);

ProductNode_POSIT11969: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT11969weight,ProductNode_POSIT1680Output_2079,ProductNode_POSIT11969Output_14815);

ProductNode_POSIT12006: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2856Output_14862,ProductNode_POSIT11969Output_14815,ProductNode_POSIT12006Output_14863);

ProductNode_POSIT12038: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2063Output_10742,ProductNode_POSIT10141Output_12553,ProductNode_POSIT12038Output_14901);

ProductNode_POSIT12070: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2069Output_10780,ProductNode_POSIT10173Output_12591,ProductNode_POSIT12070Output_14939);

SumNode_POSIT2869: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT12070Output_14939,ProductNode_POSIT12038Output_14901,SumNode_POSIT2869Output_14940);

ProductNode_POSIT12071: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2869Output_14940,ProductNode_POSIT12006Output_14863,ProductNode_POSIT12071Output_14941);

ProductNode_POSIT12073: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT12073weight,ProductNode_POSIT1784Output_2207,ProductNode_POSIT12073Output_14943);

ProductNode_POSIT12110: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2880Output_14990,ProductNode_POSIT12073Output_14943,ProductNode_POSIT12110Output_14991);

ProductNode_POSIT12142: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2087Output_10870,ProductNode_POSIT10245Output_12681,ProductNode_POSIT12142Output_15029);

ProductNode_POSIT12174: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2093Output_10908,ProductNode_POSIT10277Output_12719,ProductNode_POSIT12174Output_15067);

SumNode_POSIT2893: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT12174Output_15067,ProductNode_POSIT12142Output_15029,SumNode_POSIT2893Output_15068);

ProductNode_POSIT12175: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2893Output_15068,ProductNode_POSIT12110Output_14991,ProductNode_POSIT12175Output_15069);

SumNode_POSIT2894: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT12175Output_15069,ProductNode_POSIT12071Output_14941,SumNode_POSIT2894Output_15070);

ProductNode_POSIT12176: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb13,SumNode_POSIT2894Output_15070,ProductNode_POSIT12176Output_15071);

SumNode_POSIT2895: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT12176Output_15071,ProductNode_POSIT11967Output_14813,SumNode_POSIT2895Output_15072);

ProductNode_POSIT12177: entity work.PositMult_23_6_comb_uid2(arch)
port map(v3,SumNode_POSIT2895Output_15072,ProductNode_POSIT12177Output_15073);

ProductNode_POSIT12197: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2900Output_15097,ProductNode_POSIT2101Output_2599,ProductNode_POSIT12197Output_15098);

ProductNode_POSIT12215: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2905Output_15120,ProductNode_POSIT2119Output_2622,ProductNode_POSIT12215Output_15121);

SumNode_POSIT2906: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT12215Output_15121,ProductNode_POSIT12197Output_15098,SumNode_POSIT2906Output_15122);

ProductNode_POSIT12216: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2906Output_15122,ProductNode_POSIT11760Output_14557,ProductNode_POSIT12216Output_15123);

ProductNode_POSIT12248: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2113Output_11002,ProductNode_POSIT10560Output_13071,ProductNode_POSIT12248Output_15161);

ProductNode_POSIT12280: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2119Output_11040,ProductNode_POSIT10592Output_13109,ProductNode_POSIT12280Output_15199);

SumNode_POSIT2919: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT12280Output_15199,ProductNode_POSIT12248Output_15161,SumNode_POSIT2919Output_15200);

ProductNode_POSIT12281: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2919Output_15200,ProductNode_POSIT12216Output_15123,ProductNode_POSIT12281Output_15201);

ProductNode_POSIT12301: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2924Output_15225,ProductNode_POSIT2101Output_2599,ProductNode_POSIT12301Output_15226);

ProductNode_POSIT12319: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2929Output_15248,ProductNode_POSIT2119Output_2622,ProductNode_POSIT12319Output_15249);

SumNode_POSIT2930: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT12319Output_15249,ProductNode_POSIT12301Output_15226,SumNode_POSIT2930Output_15250);

ProductNode_POSIT12320: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2930Output_15250,ProductNode_POSIT11864Output_14685,ProductNode_POSIT12320Output_15251);

ProductNode_POSIT12352: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2137Output_11130,ProductNode_POSIT10664Output_13199,ProductNode_POSIT12352Output_15289);

ProductNode_POSIT12384: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2143Output_11168,ProductNode_POSIT10696Output_13237,ProductNode_POSIT12384Output_15327);

SumNode_POSIT2943: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT12384Output_15327,ProductNode_POSIT12352Output_15289,SumNode_POSIT2943Output_15328);

ProductNode_POSIT12385: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2943Output_15328,ProductNode_POSIT12320Output_15251,ProductNode_POSIT12385Output_15329);

SumNode_POSIT2944: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT12385Output_15329,ProductNode_POSIT12281Output_15201,SumNode_POSIT2944Output_15330);

ProductNode_POSIT12386: entity work.PositMult_23_6_comb_uid2(arch)
port map(v13,SumNode_POSIT2944Output_15330,ProductNode_POSIT12386Output_15331);

ProductNode_POSIT12425: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2955Output_15380,ProductNode_POSIT11969Output_14815,ProductNode_POSIT12425Output_15381);

ProductNode_POSIT12457: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2162Output_11260,ProductNode_POSIT10560Output_13071,ProductNode_POSIT12457Output_15419);

ProductNode_POSIT12489: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2168Output_11298,ProductNode_POSIT10592Output_13109,ProductNode_POSIT12489Output_15457);

SumNode_POSIT2968: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT12489Output_15457,ProductNode_POSIT12457Output_15419,SumNode_POSIT2968Output_15458);

ProductNode_POSIT12490: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2968Output_15458,ProductNode_POSIT12425Output_15381,ProductNode_POSIT12490Output_15459);

ProductNode_POSIT12529: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2979Output_15508,ProductNode_POSIT12073Output_14943,ProductNode_POSIT12529Output_15509);

ProductNode_POSIT12561: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2186Output_11388,ProductNode_POSIT10664Output_13199,ProductNode_POSIT12561Output_15547);

ProductNode_POSIT12593: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2192Output_11426,ProductNode_POSIT10696Output_13237,ProductNode_POSIT12593Output_15585);

SumNode_POSIT2992: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT12593Output_15585,ProductNode_POSIT12561Output_15547,SumNode_POSIT2992Output_15586);

ProductNode_POSIT12594: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2992Output_15586,ProductNode_POSIT12529Output_15509,ProductNode_POSIT12594Output_15587);

SumNode_POSIT2993: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT12594Output_15587,ProductNode_POSIT12490Output_15459,SumNode_POSIT2993Output_15588);

ProductNode_POSIT12595: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb13,SumNode_POSIT2993Output_15588,ProductNode_POSIT12595Output_15589);

SumNode_POSIT2994: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT12595Output_15589,ProductNode_POSIT12386Output_15331,SumNode_POSIT2994Output_15590);

ProductNode_POSIT12596: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb3,SumNode_POSIT2994Output_15590,ProductNode_POSIT12596Output_15591);

SumNode_POSIT2995: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT12596Output_15591,ProductNode_POSIT12177Output_15073,SumNode_POSIT2995Output_15592);

ProductNode_POSIT12597: entity work.PositMult_23_6_comb_uid2(arch)
port map(v4,SumNode_POSIT2995Output_15592,ProductNode_POSIT12597Output_15593);

ProductNode_POSIT12599: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT12599weight,ProductNode_POSIT2519Output_3117,ProductNode_POSIT12599Output_15595);

ProductNode_POSIT12608: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2997Output_15605,ProductNode_POSIT5883Output_7281,ProductNode_POSIT12608Output_15606);

ProductNode_POSIT12616: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2999Output_15615,ProductNode_POSIT5891Output_7291,ProductNode_POSIT12616Output_15616);

SumNode_POSIT3000: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT12616Output_15616,ProductNode_POSIT12608Output_15606,SumNode_POSIT3000Output_15617);

ProductNode_POSIT12617: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT3000Output_15617,ProductNode_POSIT2521Output_3119,ProductNode_POSIT12617Output_15618);

ProductNode_POSIT12626: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT3002Output_15628,ProductNode_POSIT5883Output_7281,ProductNode_POSIT12626Output_15629);

ProductNode_POSIT12634: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT3004Output_15638,ProductNode_POSIT5891Output_7291,ProductNode_POSIT12634Output_15639);

SumNode_POSIT3005: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT12634Output_15639,ProductNode_POSIT12626Output_15629,SumNode_POSIT3005Output_15640);

ProductNode_POSIT12635: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT3005Output_15640,ProductNode_POSIT2539Output_3142,ProductNode_POSIT12635Output_15641);

SumNode_POSIT3006: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT12635Output_15641,ProductNode_POSIT12617Output_15618,SumNode_POSIT3006Output_15642);

ProductNode_POSIT12636: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT3006Output_15642,ProductNode_POSIT12599Output_15595,ProductNode_POSIT12636Output_15643);

ProductNode_POSIT12668: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2213Output_11522,ProductNode_POSIT10980Output_13591,ProductNode_POSIT12668Output_15681);

ProductNode_POSIT12700: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2219Output_11560,ProductNode_POSIT11012Output_13629,ProductNode_POSIT12700Output_15719);

SumNode_POSIT3019: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT12700Output_15719,ProductNode_POSIT12668Output_15681,SumNode_POSIT3019Output_15720);

ProductNode_POSIT12701: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT3019Output_15720,ProductNode_POSIT12636Output_15643,ProductNode_POSIT12701Output_15721);

ProductNode_POSIT12703: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT12703weight,ProductNode_POSIT2623Output_3245,ProductNode_POSIT12703Output_15723);

ProductNode_POSIT12712: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT3021Output_15733,ProductNode_POSIT5883Output_7281,ProductNode_POSIT12712Output_15734);

ProductNode_POSIT12720: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT3023Output_15743,ProductNode_POSIT5891Output_7291,ProductNode_POSIT12720Output_15744);

SumNode_POSIT3024: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT12720Output_15744,ProductNode_POSIT12712Output_15734,SumNode_POSIT3024Output_15745);

ProductNode_POSIT12721: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT3024Output_15745,ProductNode_POSIT2521Output_3119,ProductNode_POSIT12721Output_15746);

ProductNode_POSIT12730: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT3026Output_15756,ProductNode_POSIT5883Output_7281,ProductNode_POSIT12730Output_15757);

ProductNode_POSIT12738: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT3028Output_15766,ProductNode_POSIT5891Output_7291,ProductNode_POSIT12738Output_15767);

SumNode_POSIT3029: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT12738Output_15767,ProductNode_POSIT12730Output_15757,SumNode_POSIT3029Output_15768);

ProductNode_POSIT12739: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT3029Output_15768,ProductNode_POSIT2539Output_3142,ProductNode_POSIT12739Output_15769);

SumNode_POSIT3030: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT12739Output_15769,ProductNode_POSIT12721Output_15746,SumNode_POSIT3030Output_15770);

ProductNode_POSIT12740: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT3030Output_15770,ProductNode_POSIT12703Output_15723,ProductNode_POSIT12740Output_15771);

ProductNode_POSIT12772: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2237Output_11650,ProductNode_POSIT11084Output_13719,ProductNode_POSIT12772Output_15809);

ProductNode_POSIT12804: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2243Output_11688,ProductNode_POSIT11116Output_13757,ProductNode_POSIT12804Output_15847);

SumNode_POSIT3043: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT12804Output_15847,ProductNode_POSIT12772Output_15809,SumNode_POSIT3043Output_15848);

ProductNode_POSIT12805: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT3043Output_15848,ProductNode_POSIT12740Output_15771,ProductNode_POSIT12805Output_15849);

SumNode_POSIT3044: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT12805Output_15849,ProductNode_POSIT12701Output_15721,SumNode_POSIT3044Output_15850);

ProductNode_POSIT12806: entity work.PositMult_23_6_comb_uid2(arch)
port map(v13,SumNode_POSIT3044Output_15850,ProductNode_POSIT12806Output_15851);

ProductNode_POSIT12808: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT12808weight,ProductNode_POSIT2519Output_3117,ProductNode_POSIT12808Output_15853);

ProductNode_POSIT12845: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT3055Output_15900,ProductNode_POSIT12808Output_15853,ProductNode_POSIT12845Output_15901);

ProductNode_POSIT12877: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2262Output_11780,ProductNode_POSIT10980Output_13591,ProductNode_POSIT12877Output_15939);

ProductNode_POSIT12909: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2268Output_11818,ProductNode_POSIT11012Output_13629,ProductNode_POSIT12909Output_15977);

SumNode_POSIT3068: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT12909Output_15977,ProductNode_POSIT12877Output_15939,SumNode_POSIT3068Output_15978);

ProductNode_POSIT12910: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT3068Output_15978,ProductNode_POSIT12845Output_15901,ProductNode_POSIT12910Output_15979);

ProductNode_POSIT12912: entity work.PositMult_23_6_comb_uid2(arch)
port map(ProductNode_POSIT12912weight,ProductNode_POSIT2623Output_3245,ProductNode_POSIT12912Output_15981);

ProductNode_POSIT12949: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT3079Output_16028,ProductNode_POSIT12912Output_15981,ProductNode_POSIT12949Output_16029);

ProductNode_POSIT12981: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2286Output_11908,ProductNode_POSIT11084Output_13719,ProductNode_POSIT12981Output_16067);

ProductNode_POSIT13013: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2292Output_11946,ProductNode_POSIT11116Output_13757,ProductNode_POSIT13013Output_16105);

SumNode_POSIT3092: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT13013Output_16105,ProductNode_POSIT12981Output_16067,SumNode_POSIT3092Output_16106);

ProductNode_POSIT13014: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT3092Output_16106,ProductNode_POSIT12949Output_16029,ProductNode_POSIT13014Output_16107);

SumNode_POSIT3093: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT13014Output_16107,ProductNode_POSIT12910Output_15979,SumNode_POSIT3093Output_16108);

ProductNode_POSIT13015: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb13,SumNode_POSIT3093Output_16108,ProductNode_POSIT13015Output_16109);

SumNode_POSIT3094: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT13015Output_16109,ProductNode_POSIT12806Output_15851,SumNode_POSIT3094Output_16110);

ProductNode_POSIT13016: entity work.PositMult_23_6_comb_uid2(arch)
port map(v3,SumNode_POSIT3094Output_16110,ProductNode_POSIT13016Output_16111);

ProductNode_POSIT13036: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT3099Output_16135,ProductNode_POSIT2940Output_3637,ProductNode_POSIT13036Output_16136);

ProductNode_POSIT13054: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT3104Output_16158,ProductNode_POSIT2958Output_3660,ProductNode_POSIT13054Output_16159);

SumNode_POSIT3105: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT13054Output_16159,ProductNode_POSIT13036Output_16136,SumNode_POSIT3105Output_16160);

ProductNode_POSIT13055: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT3105Output_16160,ProductNode_POSIT12599Output_15595,ProductNode_POSIT13055Output_16161);

ProductNode_POSIT13087: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2312Output_12040,ProductNode_POSIT11399Output_14109,ProductNode_POSIT13087Output_16199);

ProductNode_POSIT13119: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2318Output_12078,ProductNode_POSIT11431Output_14147,ProductNode_POSIT13119Output_16237);

SumNode_POSIT3118: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT13119Output_16237,ProductNode_POSIT13087Output_16199,SumNode_POSIT3118Output_16238);

ProductNode_POSIT13120: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT3118Output_16238,ProductNode_POSIT13055Output_16161,ProductNode_POSIT13120Output_16239);

ProductNode_POSIT13140: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT3123Output_16263,ProductNode_POSIT2940Output_3637,ProductNode_POSIT13140Output_16264);

ProductNode_POSIT13158: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT3128Output_16286,ProductNode_POSIT2958Output_3660,ProductNode_POSIT13158Output_16287);

SumNode_POSIT3129: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT13158Output_16287,ProductNode_POSIT13140Output_16264,SumNode_POSIT3129Output_16288);

ProductNode_POSIT13159: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT3129Output_16288,ProductNode_POSIT12703Output_15723,ProductNode_POSIT13159Output_16289);

ProductNode_POSIT13191: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2336Output_12168,ProductNode_POSIT11503Output_14237,ProductNode_POSIT13191Output_16327);

ProductNode_POSIT13223: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2342Output_12206,ProductNode_POSIT11535Output_14275,ProductNode_POSIT13223Output_16365);

SumNode_POSIT3142: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT13223Output_16365,ProductNode_POSIT13191Output_16327,SumNode_POSIT3142Output_16366);

ProductNode_POSIT13224: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT3142Output_16366,ProductNode_POSIT13159Output_16289,ProductNode_POSIT13224Output_16367);

SumNode_POSIT3143: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT13224Output_16367,ProductNode_POSIT13120Output_16239,SumNode_POSIT3143Output_16368);

ProductNode_POSIT13225: entity work.PositMult_23_6_comb_uid2(arch)
port map(v13,SumNode_POSIT3143Output_16368,ProductNode_POSIT13225Output_16369);

ProductNode_POSIT13264: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT3154Output_16418,ProductNode_POSIT12808Output_15853,ProductNode_POSIT13264Output_16419);

ProductNode_POSIT13296: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2361Output_12298,ProductNode_POSIT11399Output_14109,ProductNode_POSIT13296Output_16457);

ProductNode_POSIT13328: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2367Output_12336,ProductNode_POSIT11431Output_14147,ProductNode_POSIT13328Output_16495);

SumNode_POSIT3167: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT13328Output_16495,ProductNode_POSIT13296Output_16457,SumNode_POSIT3167Output_16496);

ProductNode_POSIT13329: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT3167Output_16496,ProductNode_POSIT13264Output_16419,ProductNode_POSIT13329Output_16497);

ProductNode_POSIT13368: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT3178Output_16546,ProductNode_POSIT12912Output_15981,ProductNode_POSIT13368Output_16547);

ProductNode_POSIT13400: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2385Output_12426,ProductNode_POSIT11503Output_14237,ProductNode_POSIT13400Output_16585);

ProductNode_POSIT13432: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT2391Output_12464,ProductNode_POSIT11535Output_14275,ProductNode_POSIT13432Output_16623);

SumNode_POSIT3191: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT13432Output_16623,ProductNode_POSIT13400Output_16585,SumNode_POSIT3191Output_16624);

ProductNode_POSIT13433: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT3191Output_16624,ProductNode_POSIT13368Output_16547,ProductNode_POSIT13433Output_16625);

SumNode_POSIT3192: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT13433Output_16625,ProductNode_POSIT13329Output_16497,SumNode_POSIT3192Output_16626);

ProductNode_POSIT13434: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb13,SumNode_POSIT3192Output_16626,ProductNode_POSIT13434Output_16627);

SumNode_POSIT3193: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT13434Output_16627,ProductNode_POSIT13225Output_16369,SumNode_POSIT3193Output_16628);

ProductNode_POSIT13435: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb3,SumNode_POSIT3193Output_16628,ProductNode_POSIT13435Output_16629);

SumNode_POSIT3194: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT13435Output_16629,ProductNode_POSIT13016Output_16111,SumNode_POSIT3194Output_16630);

ProductNode_POSIT13436: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb4,SumNode_POSIT3194Output_16630,ProductNode_POSIT13436Output_16631);

SumNode_POSIT3195: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT13436Output_16631,ProductNode_POSIT12597Output_15593,SumNode_POSIT3195Output_16632);

ProductNode_POSIT13437: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb12,SumNode_POSIT3195Output_16632,ProductNode_POSIT13437Output_16633);

SumNode_POSIT3196: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT13437Output_16633,ProductNode_POSIT11758Output_14555,SumNode_POSIT3196Output_16634);

ProductNode_POSIT13438: entity work.PositMult_23_6_comb_uid2(arch)
port map(vb6,SumNode_POSIT3196Output_16634,ProductNode_POSIT13438Output_16635);

SumNode_POSIT3197: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT13438Output_16635,ProductNode_POSIT10079Output_12477,SumNode_POSIT3197Output_16636);

ProductNode_POSIT13439: entity work.PositMult_23_6_comb_uid2(arch)
port map(SumNode_POSIT3197Output_16636,ProductNode_POSIT6720Output_8319,ProductNode_POSIT13439Output_16637);

SumNode_POSIT3198: entity work.PositAdd_23_6_F0_uid2(arch)
port map(ProductNode_POSIT13439Output_16637,ProductNode_POSIT6719Output_8318,SumNode_POSIT3198Output_16638);

vout <= SumNode_POSIT3198Output_16638;
 
end architecture;

--------------------------------------------------------------------------------
--                    SmallMultTableP3x3r6XuYu_comb_uid33
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2007-2012)
--------------------------------------------------------------------------------
library ieee; 
use ieee.std_logic_1164.all;
library work;
entity SmallMultTableP3x3r6XuYu_comb_uid33 is
   port ( X : in  std_logic_vector(5 downto 0);
          Y : out  std_logic_vector(5 downto 0)   );
end entity;

architecture arch of SmallMultTableP3x3r6XuYu_comb_uid33 is
signal TableOut :  std_logic_vector(5 downto 0);
begin
  with X select TableOut <= 
   "000000" when "000000",
   "000000" when "000001",
   "000000" when "000010",
   "000000" when "000011",
   "000000" when "000100",
   "000000" when "000101",
   "000000" when "000110",
   "000000" when "000111",
   "000000" when "001000",
   "000001" when "001001",
   "000010" when "001010",
   "000011" when "001011",
   "000100" when "001100",
   "000101" when "001101",
   "000110" when "001110",
   "000111" when "001111",
   "000000" when "010000",
   "000010" when "010001",
   "000100" when "010010",
   "000110" when "010011",
   "001000" when "010100",
   "001010" when "010101",
   "001100" when "010110",
   "001110" when "010111",
   "000000" when "011000",
   "000011" when "011001",
   "000110" when "011010",
   "001001" when "011011",
   "001100" when "011100",
   "001111" when "011101",
   "010010" when "011110",
   "010101" when "011111",
   "000000" when "100000",
   "000100" when "100001",
   "001000" when "100010",
   "001100" when "100011",
   "010000" when "100100",
   "010100" when "100101",
   "011000" when "100110",
   "011100" when "100111",
   "000000" when "101000",
   "000101" when "101001",
   "001010" when "101010",
   "001111" when "101011",
   "010100" when "101100",
   "011001" when "101101",
   "011110" when "101110",
   "100011" when "101111",
   "000000" when "110000",
   "000110" when "110001",
   "001100" when "110010",
   "010010" when "110011",
   "011000" when "110100",
   "011110" when "110101",
   "100100" when "110110",
   "101010" when "110111",
   "000000" when "111000",
   "000111" when "111001",
   "001110" when "111010",
   "010101" when "111011",
   "011100" when "111100",
   "100011" when "111101",
   "101010" when "111110",
   "110001" when "111111",
   "------" when others;
    Y <= TableOut;
end architecture;

--------------------------------------------------------------------------------
--                    SmallMultTableP3x3r6XuYu_comb_uid68
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2007-2012)
--------------------------------------------------------------------------------
library ieee; 
use ieee.std_logic_1164.all;
library work;
entity SmallMultTableP3x3r6XuYu_comb_uid68 is
   port ( X : in  std_logic_vector(5 downto 0);
          Y : out  std_logic_vector(5 downto 0)   );
end entity;

architecture arch of SmallMultTableP3x3r6XuYu_comb_uid68 is
signal TableOut :  std_logic_vector(5 downto 0);
begin
  with X select TableOut <= 
   "000000" when "000000",
   "000000" when "000001",
   "000000" when "000010",
   "000000" when "000011",
   "000000" when "000100",
   "000000" when "000101",
   "000000" when "000110",
   "000000" when "000111",
   "000000" when "001000",
   "000001" when "001001",
   "000010" when "001010",
   "000011" when "001011",
   "000100" when "001100",
   "000101" when "001101",
   "000110" when "001110",
   "000111" when "001111",
   "000000" when "010000",
   "000010" when "010001",
   "000100" when "010010",
   "000110" when "010011",
   "001000" when "010100",
   "001010" when "010101",
   "001100" when "010110",
   "001110" when "010111",
   "000000" when "011000",
   "000011" when "011001",
   "000110" when "011010",
   "001001" when "011011",
   "001100" when "011100",
   "001111" when "011101",
   "010010" when "011110",
   "010101" when "011111",
   "000000" when "100000",
   "000100" when "100001",
   "001000" when "100010",
   "001100" when "100011",
   "010000" when "100100",
   "010100" when "100101",
   "011000" when "100110",
   "011100" when "100111",
   "000000" when "101000",
   "000101" when "101001",
   "001010" when "101010",
   "001111" when "101011",
   "010100" when "101100",
   "011001" when "101101",
   "011110" when "101110",
   "100011" when "101111",
   "000000" when "110000",
   "000110" when "110001",
   "001100" when "110010",
   "010010" when "110011",
   "011000" when "110100",
   "011110" when "110101",
   "100100" when "110110",
   "101010" when "110111",
   "000000" when "111000",
   "000111" when "111001",
   "001110" when "111010",
   "010101" when "111011",
   "011100" when "111100",
   "100011" when "111101",
   "101010" when "111110",
   "110001" when "111111",
   "------" when others;
    Y <= TableOut;
end architecture;

--------------------------------------------------------------------------------
--                    SmallMultTableP3x3r6XuYu_comb_uid103
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2007-2012)
--------------------------------------------------------------------------------
library ieee; 
use ieee.std_logic_1164.all;
library work;
entity SmallMultTableP3x3r6XuYu_comb_uid103 is
   port ( X : in  std_logic_vector(5 downto 0);
          Y : out  std_logic_vector(5 downto 0)   );
end entity;

architecture arch of SmallMultTableP3x3r6XuYu_comb_uid103 is
signal TableOut :  std_logic_vector(5 downto 0);
begin
  with X select TableOut <= 
   "000000" when "000000",
   "000000" when "000001",
   "000000" when "000010",
   "000000" when "000011",
   "000000" when "000100",
   "000000" when "000101",
   "000000" when "000110",
   "000000" when "000111",
   "000000" when "001000",
   "000001" when "001001",
   "000010" when "001010",
   "000011" when "001011",
   "000100" when "001100",
   "000101" when "001101",
   "000110" when "001110",
   "000111" when "001111",
   "000000" when "010000",
   "000010" when "010001",
   "000100" when "010010",
   "000110" when "010011",
   "001000" when "010100",
   "001010" when "010101",
   "001100" when "010110",
   "001110" when "010111",
   "000000" when "011000",
   "000011" when "011001",
   "000110" when "011010",
   "001001" when "011011",
   "001100" when "011100",
   "001111" when "011101",
   "010010" when "011110",
   "010101" when "011111",
   "000000" when "100000",
   "000100" when "100001",
   "001000" when "100010",
   "001100" when "100011",
   "010000" when "100100",
   "010100" when "100101",
   "011000" when "100110",
   "011100" when "100111",
   "000000" when "101000",
   "000101" when "101001",
   "001010" when "101010",
   "001111" when "101011",
   "010100" when "101100",
   "011001" when "101101",
   "011110" when "101110",
   "100011" when "101111",
   "000000" when "110000",
   "000110" when "110001",
   "001100" when "110010",
   "010010" when "110011",
   "011000" when "110100",
   "011110" when "110101",
   "100100" when "110110",
   "101010" when "110111",
   "000000" when "111000",
   "000111" when "111001",
   "001110" when "111010",
   "010101" when "111011",
   "011100" when "111100",
   "100011" when "111101",
   "101010" when "111110",
   "110001" when "111111",
   "------" when others;
    Y <= TableOut;
end architecture;

--------------------------------------------------------------------------------
--                    SmallMultTableP3x3r6XuYu_comb_uid138
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2007-2012)
--------------------------------------------------------------------------------
library ieee; 
use ieee.std_logic_1164.all;
library work;
entity SmallMultTableP3x3r6XuYu_comb_uid138 is
   port ( X : in  std_logic_vector(5 downto 0);
          Y : out  std_logic_vector(5 downto 0)   );
end entity;

architecture arch of SmallMultTableP3x3r6XuYu_comb_uid138 is
signal TableOut :  std_logic_vector(5 downto 0);
begin
  with X select TableOut <= 
   "000000" when "000000",
   "000000" when "000001",
   "000000" when "000010",
   "000000" when "000011",
   "000000" when "000100",
   "000000" when "000101",
   "000000" when "000110",
   "000000" when "000111",
   "000000" when "001000",
   "000001" when "001001",
   "000010" when "001010",
   "000011" when "001011",
   "000100" when "001100",
   "000101" when "001101",
   "000110" when "001110",
   "000111" when "001111",
   "000000" when "010000",
   "000010" when "010001",
   "000100" when "010010",
   "000110" when "010011",
   "001000" when "010100",
   "001010" when "010101",
   "001100" when "010110",
   "001110" when "010111",
   "000000" when "011000",
   "000011" when "011001",
   "000110" when "011010",
   "001001" when "011011",
   "001100" when "011100",
   "001111" when "011101",
   "010010" when "011110",
   "010101" when "011111",
   "000000" when "100000",
   "000100" when "100001",
   "001000" when "100010",
   "001100" when "100011",
   "010000" when "100100",
   "010100" when "100101",
   "011000" when "100110",
   "011100" when "100111",
   "000000" when "101000",
   "000101" when "101001",
   "001010" when "101010",
   "001111" when "101011",
   "010100" when "101100",
   "011001" when "101101",
   "011110" when "101110",
   "100011" when "101111",
   "000000" when "110000",
   "000110" when "110001",
   "001100" when "110010",
   "010010" when "110011",
   "011000" when "110100",
   "011110" when "110101",
   "100100" when "110110",
   "101010" when "110111",
   "000000" when "111000",
   "000111" when "111001",
   "001110" when "111010",
   "010101" when "111011",
   "011100" when "111100",
   "100011" when "111101",
   "101010" when "111110",
   "110001" when "111111",
   "------" when others;
    Y <= TableOut;
end architecture;

--------------------------------------------------------------------------------
--                               Compressor_6_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Popa, Illyes Kinga, 2012
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_6_3 is
   port ( X0 : in  std_logic_vector(5 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_6_3 is
signal X :  std_logic_vector(5 downto 0);
begin
   X <=X0 ;
   with X select R <= 
      "000" when "000000", 
      "001" when "000001", 
      "001" when "000010", 
      "010" when "000011", 
      "001" when "000100", 
      "010" when "000101", 
      "010" when "000110", 
      "011" when "000111", 
      "001" when "001000", 
      "010" when "001001", 
      "010" when "001010", 
      "011" when "001011", 
      "010" when "001100", 
      "011" when "001101", 
      "011" when "001110", 
      "100" when "001111", 
      "001" when "010000", 
      "010" when "010001", 
      "010" when "010010", 
      "011" when "010011", 
      "010" when "010100", 
      "011" when "010101", 
      "011" when "010110", 
      "100" when "010111", 
      "010" when "011000", 
      "011" when "011001", 
      "011" when "011010", 
      "100" when "011011", 
      "011" when "011100", 
      "100" when "011101", 
      "100" when "011110", 
      "101" when "011111", 
      "001" when "100000", 
      "010" when "100001", 
      "010" when "100010", 
      "011" when "100011", 
      "010" when "100100", 
      "011" when "100101", 
      "011" when "100110", 
      "100" when "100111", 
      "010" when "101000", 
      "011" when "101001", 
      "011" when "101010", 
      "100" when "101011", 
      "011" when "101100", 
      "100" when "101101", 
      "100" when "101110", 
      "101" when "101111", 
      "010" when "110000", 
      "011" when "110001", 
      "011" when "110010", 
      "100" when "110011", 
      "011" when "110100", 
      "100" when "110101", 
      "100" when "110110", 
      "101" when "110111", 
      "011" when "111000", 
      "100" when "111001", 
      "100" when "111010", 
      "101" when "111011", 
      "100" when "111100", 
      "101" when "111101", 
      "101" when "111110", 
      "110" when "111111", 
      "---" when others;

end architecture;

--------------------------------------------------------------------------------
--                              Compressor_14_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Popa, Illyes Kinga, 2012
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_14_3 is
   port ( X0 : in  std_logic_vector(3 downto 0);
          X1 : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_14_3 is
signal X :  std_logic_vector(4 downto 0);
begin
   X <=X1 & X0 ;
   with X select R <= 
      "000" when "00000", 
      "001" when "00001", 
      "001" when "00010", 
      "010" when "00011", 
      "001" when "00100", 
      "010" when "00101", 
      "010" when "00110", 
      "011" when "00111", 
      "001" when "01000", 
      "010" when "01001", 
      "010" when "01010", 
      "011" when "01011", 
      "010" when "01100", 
      "011" when "01101", 
      "011" when "01110", 
      "100" when "01111", 
      "010" when "10000", 
      "011" when "10001", 
      "011" when "10010", 
      "100" when "10011", 
      "011" when "10100", 
      "100" when "10101", 
      "100" when "10110", 
      "101" when "10111", 
      "011" when "11000", 
      "100" when "11001", 
      "100" when "11010", 
      "101" when "11011", 
      "100" when "11100", 
      "101" when "11101", 
      "101" when "11110", 
      "110" when "11111", 
      "---" when others;

end architecture;

--------------------------------------------------------------------------------
--                               Compressor_5_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Popa, Illyes Kinga, 2012
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_5_3 is
   port ( X0 : in  std_logic_vector(4 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_5_3 is
signal X :  std_logic_vector(4 downto 0);
begin
   X <=X0 ;
   with X select R <= 
      "000" when "00000", 
      "001" when "00001", 
      "001" when "00010", 
      "010" when "00011", 
      "001" when "00100", 
      "010" when "00101", 
      "010" when "00110", 
      "011" when "00111", 
      "001" when "01000", 
      "010" when "01001", 
      "010" when "01010", 
      "011" when "01011", 
      "010" when "01100", 
      "011" when "01101", 
      "011" when "01110", 
      "100" when "01111", 
      "001" when "10000", 
      "010" when "10001", 
      "010" when "10010", 
      "011" when "10011", 
      "010" when "10100", 
      "011" when "10101", 
      "011" when "10110", 
      "100" when "10111", 
      "010" when "11000", 
      "011" when "11001", 
      "011" when "11010", 
      "100" when "11011", 
      "011" when "11100", 
      "100" when "11101", 
      "100" when "11110", 
      "101" when "11111", 
      "---" when others;

end architecture;

--------------------------------------------------------------------------------
--                               Compressor_4_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Popa, Illyes Kinga, 2012
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_4_3 is
   port ( X0 : in  std_logic_vector(3 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_4_3 is
signal X :  std_logic_vector(3 downto 0);
begin
   X <=X0 ;
   with X select R <= 
      "000" when "0000", 
      "001" when "0001", 
      "001" when "0010", 
      "010" when "0011", 
      "001" when "0100", 
      "010" when "0101", 
      "010" when "0110", 
      "011" when "0111", 
      "001" when "1000", 
      "010" when "1001", 
      "010" when "1010", 
      "011" when "1011", 
      "010" when "1100", 
      "011" when "1101", 
      "011" when "1110", 
      "100" when "1111", 
      "---" when others;

end architecture;

--------------------------------------------------------------------------------
--                              Compressor_23_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Popa, Illyes Kinga, 2012
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_23_3 is
   port ( X0 : in  std_logic_vector(2 downto 0);
          X1 : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_23_3 is
signal X :  std_logic_vector(4 downto 0);
begin
   X <=X1 & X0 ;
   with X select R <= 
      "000" when "00000", 
      "001" when "00001", 
      "001" when "00010", 
      "010" when "00011", 
      "001" when "00100", 
      "010" when "00101", 
      "010" when "00110", 
      "011" when "00111", 
      "010" when "01000", 
      "011" when "01001", 
      "011" when "01010", 
      "100" when "01011", 
      "011" when "01100", 
      "100" when "01101", 
      "100" when "01110", 
      "101" when "01111", 
      "010" when "10000", 
      "011" when "10001", 
      "011" when "10010", 
      "100" when "10011", 
      "011" when "10100", 
      "100" when "10101", 
      "100" when "10110", 
      "101" when "10111", 
      "100" when "11000", 
      "101" when "11001", 
      "101" when "11010", 
      "110" when "11011", 
      "101" when "11100", 
      "110" when "11101", 
      "110" when "11110", 
      "111" when "11111", 
      "---" when others;

end architecture;

--------------------------------------------------------------------------------
--                              Compressor_13_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Popa, Illyes Kinga, 2012
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_13_3 is
   port ( X0 : in  std_logic_vector(2 downto 0);
          X1 : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_13_3 is
signal X :  std_logic_vector(3 downto 0);
begin
   X <=X1 & X0 ;
   with X select R <= 
      "000" when "0000", 
      "001" when "0001", 
      "001" when "0010", 
      "010" when "0011", 
      "001" when "0100", 
      "010" when "0101", 
      "010" when "0110", 
      "011" when "0111", 
      "010" when "1000", 
      "011" when "1001", 
      "011" when "1010", 
      "100" when "1011", 
      "011" when "1100", 
      "100" when "1101", 
      "100" when "1110", 
      "101" when "1111", 
      "---" when others;

end architecture;

--------------------------------------------------------------------------------
--                               Compressor_3_2
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Popa, Illyes Kinga, 2012
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_3_2 is
   port ( X0 : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of Compressor_3_2 is
signal X :  std_logic_vector(2 downto 0);
begin
   X <=X0 ;
   with X select R <= 
      "00" when "000", 
      "01" when "001", 
      "01" when "010", 
      "10" when "011", 
      "01" when "100", 
      "10" when "101", 
      "10" when "110", 
      "11" when "111", 
      "--" when others;

end architecture;

--------------------------------------------------------------------------------
--                             LZOC_99_comb_uid6
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007)
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LZOC_99_comb_uid6 is
   port ( I : in  std_logic_vector(98 downto 0);
          OZB : in  std_logic;
          O : out  std_logic_vector(6 downto 0)   );
end entity;

architecture arch of LZOC_99_comb_uid6 is
signal sozb :  std_logic;
signal level7 :  std_logic_vector(127 downto 0);
signal digit7 :  std_logic;
signal level6 :  std_logic_vector(63 downto 0);
signal digit6 :  std_logic;
signal level5 :  std_logic_vector(31 downto 0);
signal digit5 :  std_logic;
signal level4 :  std_logic_vector(15 downto 0);
signal digit4 :  std_logic;
signal level3 :  std_logic_vector(7 downto 0);
signal digit3 :  std_logic;
signal level2 :  std_logic_vector(3 downto 0);
signal digit2 :  std_logic;
signal level1 :  std_logic_vector(1 downto 0);
signal digit1 :  std_logic;
begin
   sozb <= OZB;
   level7<= I& (28 downto 0 => not(sozb));
   digit7<= '1' when level7(127 downto 64) = (127 downto 64 => sozb) else '0';
   level6<= level7(63 downto 0) when digit7='1' else level7(127 downto 64);
   digit6<= '1' when level6(63 downto 32) = (63 downto 32 => sozb) else '0';
   level5<= level6(31 downto 0) when digit6='1' else level6(63 downto 32);
   digit5<= '1' when level5(31 downto 16) = (31 downto 16 => sozb) else '0';
   level4<= level5(15 downto 0) when digit5='1' else level5(31 downto 16);
   digit4<= '1' when level4(15 downto 8) = (15 downto 8 => sozb) else '0';
   level3<= level4(7 downto 0) when digit4='1' else level4(15 downto 8);
   digit3<= '1' when level3(7 downto 4) = (7 downto 4 => sozb) else '0';
   level2<= level3(3 downto 0) when digit3='1' else level3(7 downto 4);
   digit2<= '1' when level2(3 downto 2) = (3 downto 2 => sozb) else '0';
   level1<= level2(1 downto 0) when digit2='1' else level2(3 downto 2);
   digit1<= '1' when level1(1 downto 1) = (1 downto 1 => sozb) else '0';
   O <= digit7 & digit6 & digit5 & digit4 & digit3 & digit2 & digit1;
end architecture;

--------------------------------------------------------------------------------
--                    LeftShifter_99_by_max_99_comb_uid10
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2011)
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LeftShifter_99_by_max_99_comb_uid10 is
   port ( X : in  std_logic_vector(98 downto 0);
          S : in  std_logic_vector(6 downto 0);
          R : out  std_logic_vector(197 downto 0)   );
end entity;

architecture arch of LeftShifter_99_by_max_99_comb_uid10 is
signal level0 :  std_logic_vector(98 downto 0);
signal ps :  std_logic_vector(6 downto 0);
signal level1 :  std_logic_vector(99 downto 0);
signal level2 :  std_logic_vector(101 downto 0);
signal level3 :  std_logic_vector(105 downto 0);
signal level4 :  std_logic_vector(113 downto 0);
signal level5 :  std_logic_vector(129 downto 0);
signal level6 :  std_logic_vector(161 downto 0);
signal level7 :  std_logic_vector(225 downto 0);
begin
   level0<= X;
   ps<= S;
   level1<= level0 & (0 downto 0 => '0') when ps(0)= '1' else     (0 downto 0 => '0') & level0;
   level2<= level1 & (1 downto 0 => '0') when ps(1)= '1' else     (1 downto 0 => '0') & level1;
   level3<= level2 & (3 downto 0 => '0') when ps(2)= '1' else     (3 downto 0 => '0') & level2;
   level4<= level3 & (7 downto 0 => '0') when ps(3)= '1' else     (7 downto 0 => '0') & level3;
   level5<= level4 & (15 downto 0 => '0') when ps(4)= '1' else     (15 downto 0 => '0') & level4;
   level6<= level5 & (31 downto 0 => '0') when ps(5)= '1' else     (31 downto 0 => '0') & level5;
   level7<= level6 & (63 downto 0 => '0') when ps(6)= '1' else     (63 downto 0 => '0') & level6;
   R <= level7(197 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                        PositDecoder_100_8_comb_uid4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Raul Murillo, 2019
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity PositDecoder_100_8_comb_uid4 is
   port ( Input : in  std_logic_vector(99 downto 0);
          Sign : out  std_logic;
          Reg : out  std_logic_vector(7 downto 0);
          Exp : out  std_logic_vector(7 downto 0);
          Frac : out  std_logic_vector(89 downto 0);
          z : out  std_logic;
          inf : out  std_logic   );
end entity;

architecture arch of PositDecoder_100_8_comb_uid4 is
   component LZOC_99_comb_uid6 is
      port ( I : in  std_logic_vector(98 downto 0);
             OZB : in  std_logic;
             O : out  std_logic_vector(6 downto 0)   );
   end component;

   component LeftShifter_99_by_max_99_comb_uid10 is
      port ( X : in  std_logic_vector(98 downto 0);
             S : in  std_logic_vector(6 downto 0);
             R : out  std_logic_vector(197 downto 0)   );
   end component;

signal nzero :  std_logic;
signal my_sign :  std_logic;
signal rep_sign :  std_logic_vector(98 downto 0);
signal twos :  std_logic_vector(98 downto 0);
signal rc :  std_logic;
signal rep_rc :  std_logic_vector(98 downto 0);
signal inv :  std_logic_vector(98 downto 0);
signal zero_var :  std_logic;
signal zc :  std_logic_vector(6 downto 0);
signal zc_sub :  std_logic_vector(6 downto 0);
signal shifted_twos :  std_logic_vector(197 downto 0);
signal tmp :  std_logic_vector(96 downto 0);
begin
-------------------------------- Special Cases --------------------------------
   nzero <= '0' when Input(98 downto 0) = 0 else '1';
   -- 1 if Input is zero
   z <= Input(99) NOR nzero;
   -- 1 if Input is infinity
   inf <= Input(99) AND (NOT nzero);
------------------------------- Extract Sign bit -------------------------------
   my_sign <= Input(99);
   Sign <= my_sign;
--------------------------- 2's Complement of Input ---------------------------
   rep_sign <= (others => my_sign);
   twos <= (rep_sign XOR Input(98 downto 0)) + my_sign;
   rc <= twos(98);
------------------------ Count leading zeros of regime ------------------------
   rep_rc <= (others => rc);
   -- Invert 2's
   inv <= rep_rc XOR twos;
   zero_var <= '0';
   LZOC_Component: LZOC_99_comb_uid6
      port map ( I => inv,
                 O => zc,
                 OZB => zero_var);
----------------------------- Shift out the regime -----------------------------
   zc_sub <= zc - 1;
   LeftShifterComponent: LeftShifter_99_by_max_99_comb_uid10
      port map ( R => shifted_twos,
                 S => zc_sub,
                 X => twos);
   tmp <= shifted_twos(96 downto 0);
------------------------ Extract fraction and exponent ------------------------
   Frac <= nzero & tmp(88 downto 0);
   Exp <= tmp(96 downto 89);
-------------------------------- Select regime --------------------------------
   Reg <= '0' & zc_sub when rc = '1' else NOT('0' & zc) + 1;
end architecture;

--------------------------------------------------------------------------------
--                             LZOC_99_comb_uid18
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007)
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LZOC_99_comb_uid18 is
   port ( I : in  std_logic_vector(98 downto 0);
          OZB : in  std_logic;
          O : out  std_logic_vector(6 downto 0)   );
end entity;

architecture arch of LZOC_99_comb_uid18 is
signal sozb :  std_logic;
signal level7 :  std_logic_vector(127 downto 0);
signal digit7 :  std_logic;
signal level6 :  std_logic_vector(63 downto 0);
signal digit6 :  std_logic;
signal level5 :  std_logic_vector(31 downto 0);
signal digit5 :  std_logic;
signal level4 :  std_logic_vector(15 downto 0);
signal digit4 :  std_logic;
signal level3 :  std_logic_vector(7 downto 0);
signal digit3 :  std_logic;
signal level2 :  std_logic_vector(3 downto 0);
signal digit2 :  std_logic;
signal level1 :  std_logic_vector(1 downto 0);
signal digit1 :  std_logic;
begin
   sozb <= OZB;
   level7<= I& (28 downto 0 => not(sozb));
   digit7<= '1' when level7(127 downto 64) = (127 downto 64 => sozb) else '0';
   level6<= level7(63 downto 0) when digit7='1' else level7(127 downto 64);
   digit6<= '1' when level6(63 downto 32) = (63 downto 32 => sozb) else '0';
   level5<= level6(31 downto 0) when digit6='1' else level6(63 downto 32);
   digit5<= '1' when level5(31 downto 16) = (31 downto 16 => sozb) else '0';
   level4<= level5(15 downto 0) when digit5='1' else level5(31 downto 16);
   digit4<= '1' when level4(15 downto 8) = (15 downto 8 => sozb) else '0';
   level3<= level4(7 downto 0) when digit4='1' else level4(15 downto 8);
   digit3<= '1' when level3(7 downto 4) = (7 downto 4 => sozb) else '0';
   level2<= level3(3 downto 0) when digit3='1' else level3(7 downto 4);
   digit2<= '1' when level2(3 downto 2) = (3 downto 2 => sozb) else '0';
   level1<= level2(1 downto 0) when digit2='1' else level2(3 downto 2);
   digit1<= '1' when level1(1 downto 1) = (1 downto 1 => sozb) else '0';
   O <= digit7 & digit6 & digit5 & digit4 & digit3 & digit2 & digit1;
end architecture;

--------------------------------------------------------------------------------
--                    LeftShifter_99_by_max_99_comb_uid22
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2011)
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LeftShifter_99_by_max_99_comb_uid22 is
   port ( X : in  std_logic_vector(98 downto 0);
          S : in  std_logic_vector(6 downto 0);
          R : out  std_logic_vector(197 downto 0)   );
end entity;

architecture arch of LeftShifter_99_by_max_99_comb_uid22 is
signal level0 :  std_logic_vector(98 downto 0);
signal ps :  std_logic_vector(6 downto 0);
signal level1 :  std_logic_vector(99 downto 0);
signal level2 :  std_logic_vector(101 downto 0);
signal level3 :  std_logic_vector(105 downto 0);
signal level4 :  std_logic_vector(113 downto 0);
signal level5 :  std_logic_vector(129 downto 0);
signal level6 :  std_logic_vector(161 downto 0);
signal level7 :  std_logic_vector(225 downto 0);
begin
   level0<= X;
   ps<= S;
   level1<= level0 & (0 downto 0 => '0') when ps(0)= '1' else     (0 downto 0 => '0') & level0;
   level2<= level1 & (1 downto 0 => '0') when ps(1)= '1' else     (1 downto 0 => '0') & level1;
   level3<= level2 & (3 downto 0 => '0') when ps(2)= '1' else     (3 downto 0 => '0') & level2;
   level4<= level3 & (7 downto 0 => '0') when ps(3)= '1' else     (7 downto 0 => '0') & level3;
   level5<= level4 & (15 downto 0 => '0') when ps(4)= '1' else     (15 downto 0 => '0') & level4;
   level6<= level5 & (31 downto 0 => '0') when ps(5)= '1' else     (31 downto 0 => '0') & level5;
   level7<= level6 & (63 downto 0 => '0') when ps(6)= '1' else     (63 downto 0 => '0') & level6;
   R <= level7(197 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                       PositDecoder_100_8_comb_uid16
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Raul Murillo, 2019
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity PositDecoder_100_8_comb_uid16 is
   port ( Input : in  std_logic_vector(99 downto 0);
          Sign : out  std_logic;
          Reg : out  std_logic_vector(7 downto 0);
          Exp : out  std_logic_vector(7 downto 0);
          Frac : out  std_logic_vector(89 downto 0);
          z : out  std_logic;
          inf : out  std_logic   );
end entity;

architecture arch of PositDecoder_100_8_comb_uid16 is
   component LZOC_99_comb_uid18 is
      port ( I : in  std_logic_vector(98 downto 0);
             OZB : in  std_logic;
             O : out  std_logic_vector(6 downto 0)   );
   end component;

   component LeftShifter_99_by_max_99_comb_uid22 is
      port ( X : in  std_logic_vector(98 downto 0);
             S : in  std_logic_vector(6 downto 0);
             R : out  std_logic_vector(197 downto 0)   );
   end component;

signal nzero :  std_logic;
signal my_sign :  std_logic;
signal rep_sign :  std_logic_vector(98 downto 0);
signal twos :  std_logic_vector(98 downto 0);
signal rc :  std_logic;
signal rep_rc :  std_logic_vector(98 downto 0);
signal inv :  std_logic_vector(98 downto 0);
signal zero_var :  std_logic;
signal zc :  std_logic_vector(6 downto 0);
signal zc_sub :  std_logic_vector(6 downto 0);
signal shifted_twos :  std_logic_vector(197 downto 0);
signal tmp :  std_logic_vector(96 downto 0);
begin
-------------------------------- Special Cases --------------------------------
   nzero <= '0' when Input(98 downto 0) = 0 else '1';
   -- 1 if Input is zero
   z <= Input(99) NOR nzero;
   -- 1 if Input is infinity
   inf <= Input(99) AND (NOT nzero);
------------------------------- Extract Sign bit -------------------------------
   my_sign <= Input(99);
   Sign <= my_sign;
--------------------------- 2's Complement of Input ---------------------------
   rep_sign <= (others => my_sign);
   twos <= (rep_sign XOR Input(98 downto 0)) + my_sign;
   rc <= twos(98);
------------------------ Count leading zeros of regime ------------------------
   rep_rc <= (others => rc);
   -- Invert 2's
   inv <= rep_rc XOR twos;
   zero_var <= '0';
   LZOC_Component: LZOC_99_comb_uid18
      port map ( I => inv,
                 O => zc,
                 OZB => zero_var);
----------------------------- Shift out the regime -----------------------------
   zc_sub <= zc - 1;
   LeftShifterComponent: LeftShifter_99_by_max_99_comb_uid22
      port map ( R => shifted_twos,
                 S => zc_sub,
                 X => twos);
   tmp <= shifted_twos(96 downto 0);
------------------------ Extract fraction and exponent ------------------------
   Frac <= nzero & tmp(88 downto 0);
   Exp <= tmp(96 downto 89);
-------------------------------- Select regime --------------------------------
   Reg <= '0' & zc_sub when rc = '1' else NOT('0' & zc) + 1;
end architecture;

--------------------------------------------------------------------------------
--                         IntAdder_181_f400_uid1117
--                   (IntAdderAlternative_181_comb_uid1121)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_181_f400_uid1117 is
   port ( X : in  std_logic_vector(180 downto 0);
          Y : in  std_logic_vector(180 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(180 downto 0)   );
end entity;

architecture arch of IntAdder_181_f400_uid1117 is
begin
   --Alternative
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--            IntMultiplier_UsingDSP_90_90_180_unsigned_comb_uid28
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Kinga Illyes, Bogdan Popa, Bogdan Pasca, 2012
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity IntMultiplier_UsingDSP_90_90_180_unsigned_comb_uid28 is
   port ( X : in  std_logic_vector(89 downto 0);
          Y : in  std_logic_vector(89 downto 0);
          R : out  std_logic_vector(179 downto 0)   );
end entity;

architecture arch of IntMultiplier_UsingDSP_90_90_180_unsigned_comb_uid28 is
   component IntAdder_181_f400_uid1117 is
      port ( X : in  std_logic_vector(180 downto 0);
             Y : in  std_logic_vector(180 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(180 downto 0)   );
   end component;

   component SmallMultTableP3x3r6XuYu_comb_uid33 is
      port ( X : in  std_logic_vector(5 downto 0);
             Y : out  std_logic_vector(5 downto 0)   );
   end component;

   component SmallMultTableP3x3r6XuYu_comb_uid68 is
      port ( X : in  std_logic_vector(5 downto 0);
             Y : out  std_logic_vector(5 downto 0)   );
   end component;

   component SmallMultTableP3x3r6XuYu_comb_uid103 is
      port ( X : in  std_logic_vector(5 downto 0);
             Y : out  std_logic_vector(5 downto 0)   );
   end component;

   component SmallMultTableP3x3r6XuYu_comb_uid138 is
      port ( X : in  std_logic_vector(5 downto 0);
             Y : out  std_logic_vector(5 downto 0)   );
   end component;

   component Compressor_6_3 is
      port ( X0 : in  std_logic_vector(5 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_14_3 is
      port ( X0 : in  std_logic_vector(3 downto 0);
             X1 : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_5_3 is
      port ( X0 : in  std_logic_vector(4 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_4_3 is
      port ( X0 : in  std_logic_vector(3 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_23_3 is
      port ( X0 : in  std_logic_vector(2 downto 0);
             X1 : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_13_3 is
      port ( X0 : in  std_logic_vector(2 downto 0);
             X1 : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_3_2 is
      port ( X0 : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

signal XX_m29 :  std_logic_vector(89 downto 0);
signal YY_m29 :  std_logic_vector(89 downto 0);
signal Xp_m29b31 :  std_logic_vector(23 downto 0);
signal Yp_m29b31 :  std_logic_vector(5 downto 0);
signal x_m29b31_0 :  std_logic_vector(2 downto 0);
signal x_m29b31_1 :  std_logic_vector(2 downto 0);
signal x_m29b31_2 :  std_logic_vector(2 downto 0);
signal x_m29b31_3 :  std_logic_vector(2 downto 0);
signal x_m29b31_4 :  std_logic_vector(2 downto 0);
signal x_m29b31_5 :  std_logic_vector(2 downto 0);
signal x_m29b31_6 :  std_logic_vector(2 downto 0);
signal x_m29b31_7 :  std_logic_vector(2 downto 0);
signal y_m29b31_0 :  std_logic_vector(2 downto 0);
signal y_m29b31_1 :  std_logic_vector(2 downto 0);
signal Y0X0_31_m29 :  std_logic_vector(5 downto 0);
signal PP31X0Y0_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w66_0 :  std_logic;
signal heap_bh30_w67_0 :  std_logic;
signal heap_bh30_w68_0 :  std_logic;
signal heap_bh30_w69_0 :  std_logic;
signal heap_bh30_w70_0 :  std_logic;
signal Y0X1_31_m29 :  std_logic_vector(5 downto 0);
signal PP31X1Y0_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w69_1 :  std_logic;
signal heap_bh30_w70_1 :  std_logic;
signal heap_bh30_w71_0 :  std_logic;
signal heap_bh30_w72_0 :  std_logic;
signal heap_bh30_w73_0 :  std_logic;
signal Y0X2_31_m29 :  std_logic_vector(5 downto 0);
signal PP31X2Y0_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w72_1 :  std_logic;
signal heap_bh30_w73_1 :  std_logic;
signal heap_bh30_w74_0 :  std_logic;
signal heap_bh30_w75_0 :  std_logic;
signal heap_bh30_w76_0 :  std_logic;
signal Y0X3_31_m29 :  std_logic_vector(5 downto 0);
signal PP31X3Y0_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w75_1 :  std_logic;
signal heap_bh30_w76_1 :  std_logic;
signal heap_bh30_w77_0 :  std_logic;
signal heap_bh30_w78_0 :  std_logic;
signal heap_bh30_w79_0 :  std_logic;
signal Y0X4_31_m29 :  std_logic_vector(5 downto 0);
signal PP31X4Y0_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w78_1 :  std_logic;
signal heap_bh30_w79_1 :  std_logic;
signal heap_bh30_w80_0 :  std_logic;
signal heap_bh30_w81_0 :  std_logic;
signal heap_bh30_w82_0 :  std_logic;
signal Y0X5_31_m29 :  std_logic_vector(5 downto 0);
signal PP31X5Y0_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w81_1 :  std_logic;
signal heap_bh30_w82_1 :  std_logic;
signal heap_bh30_w83_0 :  std_logic;
signal heap_bh30_w84_0 :  std_logic;
signal heap_bh30_w85_0 :  std_logic;
signal Y0X6_31_m29 :  std_logic_vector(5 downto 0);
signal PP31X6Y0_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w84_1 :  std_logic;
signal heap_bh30_w85_1 :  std_logic;
signal heap_bh30_w86_0 :  std_logic;
signal heap_bh30_w87_0 :  std_logic;
signal heap_bh30_w88_0 :  std_logic;
signal Y0X7_31_m29 :  std_logic_vector(5 downto 0);
signal PP31X7Y0_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w87_1 :  std_logic;
signal heap_bh30_w88_1 :  std_logic;
signal heap_bh30_w89_0 :  std_logic;
signal heap_bh30_w90_0 :  std_logic;
signal heap_bh30_w91_0 :  std_logic;
signal Y1X0_31_m29 :  std_logic_vector(5 downto 0);
signal PP31X0Y1_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w68_1 :  std_logic;
signal heap_bh30_w69_2 :  std_logic;
signal heap_bh30_w70_2 :  std_logic;
signal heap_bh30_w71_1 :  std_logic;
signal heap_bh30_w72_2 :  std_logic;
signal heap_bh30_w73_2 :  std_logic;
signal Y1X1_31_m29 :  std_logic_vector(5 downto 0);
signal PP31X1Y1_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w71_2 :  std_logic;
signal heap_bh30_w72_3 :  std_logic;
signal heap_bh30_w73_3 :  std_logic;
signal heap_bh30_w74_1 :  std_logic;
signal heap_bh30_w75_2 :  std_logic;
signal heap_bh30_w76_2 :  std_logic;
signal Y1X2_31_m29 :  std_logic_vector(5 downto 0);
signal PP31X2Y1_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w74_2 :  std_logic;
signal heap_bh30_w75_3 :  std_logic;
signal heap_bh30_w76_3 :  std_logic;
signal heap_bh30_w77_1 :  std_logic;
signal heap_bh30_w78_2 :  std_logic;
signal heap_bh30_w79_2 :  std_logic;
signal Y1X3_31_m29 :  std_logic_vector(5 downto 0);
signal PP31X3Y1_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w77_2 :  std_logic;
signal heap_bh30_w78_3 :  std_logic;
signal heap_bh30_w79_3 :  std_logic;
signal heap_bh30_w80_1 :  std_logic;
signal heap_bh30_w81_2 :  std_logic;
signal heap_bh30_w82_2 :  std_logic;
signal Y1X4_31_m29 :  std_logic_vector(5 downto 0);
signal PP31X4Y1_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w80_2 :  std_logic;
signal heap_bh30_w81_3 :  std_logic;
signal heap_bh30_w82_3 :  std_logic;
signal heap_bh30_w83_1 :  std_logic;
signal heap_bh30_w84_2 :  std_logic;
signal heap_bh30_w85_2 :  std_logic;
signal Y1X5_31_m29 :  std_logic_vector(5 downto 0);
signal PP31X5Y1_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w83_2 :  std_logic;
signal heap_bh30_w84_3 :  std_logic;
signal heap_bh30_w85_3 :  std_logic;
signal heap_bh30_w86_1 :  std_logic;
signal heap_bh30_w87_2 :  std_logic;
signal heap_bh30_w88_2 :  std_logic;
signal Y1X6_31_m29 :  std_logic_vector(5 downto 0);
signal PP31X6Y1_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w86_2 :  std_logic;
signal heap_bh30_w87_3 :  std_logic;
signal heap_bh30_w88_3 :  std_logic;
signal heap_bh30_w89_1 :  std_logic;
signal heap_bh30_w90_1 :  std_logic;
signal heap_bh30_w91_1 :  std_logic;
signal Y1X7_31_m29 :  std_logic_vector(5 downto 0);
signal PP31X7Y1_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w89_2 :  std_logic;
signal heap_bh30_w90_2 :  std_logic;
signal heap_bh30_w91_2 :  std_logic;
signal heap_bh30_w92_0 :  std_logic;
signal heap_bh30_w93_0 :  std_logic;
signal heap_bh30_w94_0 :  std_logic;
signal Xp_m29b66 :  std_logic_vector(23 downto 0);
signal Yp_m29b66 :  std_logic_vector(5 downto 0);
signal x_m29b66_0 :  std_logic_vector(2 downto 0);
signal x_m29b66_1 :  std_logic_vector(2 downto 0);
signal x_m29b66_2 :  std_logic_vector(2 downto 0);
signal x_m29b66_3 :  std_logic_vector(2 downto 0);
signal x_m29b66_4 :  std_logic_vector(2 downto 0);
signal x_m29b66_5 :  std_logic_vector(2 downto 0);
signal x_m29b66_6 :  std_logic_vector(2 downto 0);
signal x_m29b66_7 :  std_logic_vector(2 downto 0);
signal y_m29b66_0 :  std_logic_vector(2 downto 0);
signal y_m29b66_1 :  std_logic_vector(2 downto 0);
signal Y0X0_66_m29 :  std_logic_vector(5 downto 0);
signal PP66X0Y0_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w42_0 :  std_logic;
signal heap_bh30_w43_0 :  std_logic;
signal heap_bh30_w44_0 :  std_logic;
signal heap_bh30_w45_0 :  std_logic;
signal heap_bh30_w46_0 :  std_logic;
signal Y0X1_66_m29 :  std_logic_vector(5 downto 0);
signal PP66X1Y0_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w45_1 :  std_logic;
signal heap_bh30_w46_1 :  std_logic;
signal heap_bh30_w47_0 :  std_logic;
signal heap_bh30_w48_0 :  std_logic;
signal heap_bh30_w49_0 :  std_logic;
signal Y0X2_66_m29 :  std_logic_vector(5 downto 0);
signal PP66X2Y0_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w48_1 :  std_logic;
signal heap_bh30_w49_1 :  std_logic;
signal heap_bh30_w50_0 :  std_logic;
signal heap_bh30_w51_0 :  std_logic;
signal heap_bh30_w52_0 :  std_logic;
signal Y0X3_66_m29 :  std_logic_vector(5 downto 0);
signal PP66X3Y0_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w51_1 :  std_logic;
signal heap_bh30_w52_1 :  std_logic;
signal heap_bh30_w53_0 :  std_logic;
signal heap_bh30_w54_0 :  std_logic;
signal heap_bh30_w55_0 :  std_logic;
signal Y0X4_66_m29 :  std_logic_vector(5 downto 0);
signal PP66X4Y0_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w54_1 :  std_logic;
signal heap_bh30_w55_1 :  std_logic;
signal heap_bh30_w56_0 :  std_logic;
signal heap_bh30_w57_0 :  std_logic;
signal heap_bh30_w58_0 :  std_logic;
signal Y0X5_66_m29 :  std_logic_vector(5 downto 0);
signal PP66X5Y0_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w57_1 :  std_logic;
signal heap_bh30_w58_1 :  std_logic;
signal heap_bh30_w59_0 :  std_logic;
signal heap_bh30_w60_0 :  std_logic;
signal heap_bh30_w61_0 :  std_logic;
signal Y0X6_66_m29 :  std_logic_vector(5 downto 0);
signal PP66X6Y0_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w60_1 :  std_logic;
signal heap_bh30_w61_1 :  std_logic;
signal heap_bh30_w62_0 :  std_logic;
signal heap_bh30_w63_0 :  std_logic;
signal heap_bh30_w64_0 :  std_logic;
signal Y0X7_66_m29 :  std_logic_vector(5 downto 0);
signal PP66X7Y0_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w63_1 :  std_logic;
signal heap_bh30_w64_1 :  std_logic;
signal heap_bh30_w65_0 :  std_logic;
signal heap_bh30_w66_1 :  std_logic;
signal heap_bh30_w67_1 :  std_logic;
signal Y1X0_66_m29 :  std_logic_vector(5 downto 0);
signal PP66X0Y1_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w44_1 :  std_logic;
signal heap_bh30_w45_2 :  std_logic;
signal heap_bh30_w46_2 :  std_logic;
signal heap_bh30_w47_1 :  std_logic;
signal heap_bh30_w48_2 :  std_logic;
signal heap_bh30_w49_2 :  std_logic;
signal Y1X1_66_m29 :  std_logic_vector(5 downto 0);
signal PP66X1Y1_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w47_2 :  std_logic;
signal heap_bh30_w48_3 :  std_logic;
signal heap_bh30_w49_3 :  std_logic;
signal heap_bh30_w50_1 :  std_logic;
signal heap_bh30_w51_2 :  std_logic;
signal heap_bh30_w52_2 :  std_logic;
signal Y1X2_66_m29 :  std_logic_vector(5 downto 0);
signal PP66X2Y1_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w50_2 :  std_logic;
signal heap_bh30_w51_3 :  std_logic;
signal heap_bh30_w52_3 :  std_logic;
signal heap_bh30_w53_1 :  std_logic;
signal heap_bh30_w54_2 :  std_logic;
signal heap_bh30_w55_2 :  std_logic;
signal Y1X3_66_m29 :  std_logic_vector(5 downto 0);
signal PP66X3Y1_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w53_2 :  std_logic;
signal heap_bh30_w54_3 :  std_logic;
signal heap_bh30_w55_3 :  std_logic;
signal heap_bh30_w56_1 :  std_logic;
signal heap_bh30_w57_2 :  std_logic;
signal heap_bh30_w58_2 :  std_logic;
signal Y1X4_66_m29 :  std_logic_vector(5 downto 0);
signal PP66X4Y1_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w56_2 :  std_logic;
signal heap_bh30_w57_3 :  std_logic;
signal heap_bh30_w58_3 :  std_logic;
signal heap_bh30_w59_1 :  std_logic;
signal heap_bh30_w60_2 :  std_logic;
signal heap_bh30_w61_2 :  std_logic;
signal Y1X5_66_m29 :  std_logic_vector(5 downto 0);
signal PP66X5Y1_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w59_2 :  std_logic;
signal heap_bh30_w60_3 :  std_logic;
signal heap_bh30_w61_3 :  std_logic;
signal heap_bh30_w62_1 :  std_logic;
signal heap_bh30_w63_2 :  std_logic;
signal heap_bh30_w64_2 :  std_logic;
signal Y1X6_66_m29 :  std_logic_vector(5 downto 0);
signal PP66X6Y1_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w62_2 :  std_logic;
signal heap_bh30_w63_3 :  std_logic;
signal heap_bh30_w64_3 :  std_logic;
signal heap_bh30_w65_1 :  std_logic;
signal heap_bh30_w66_2 :  std_logic;
signal heap_bh30_w67_2 :  std_logic;
signal Y1X7_66_m29 :  std_logic_vector(5 downto 0);
signal PP66X7Y1_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w65_2 :  std_logic;
signal heap_bh30_w66_3 :  std_logic;
signal heap_bh30_w67_3 :  std_logic;
signal heap_bh30_w68_2 :  std_logic;
signal heap_bh30_w69_3 :  std_logic;
signal heap_bh30_w70_3 :  std_logic;
signal Xp_m29b101 :  std_logic_vector(23 downto 0);
signal Yp_m29b101 :  std_logic_vector(5 downto 0);
signal x_m29b101_0 :  std_logic_vector(2 downto 0);
signal x_m29b101_1 :  std_logic_vector(2 downto 0);
signal x_m29b101_2 :  std_logic_vector(2 downto 0);
signal x_m29b101_3 :  std_logic_vector(2 downto 0);
signal x_m29b101_4 :  std_logic_vector(2 downto 0);
signal x_m29b101_5 :  std_logic_vector(2 downto 0);
signal x_m29b101_6 :  std_logic_vector(2 downto 0);
signal x_m29b101_7 :  std_logic_vector(2 downto 0);
signal y_m29b101_0 :  std_logic_vector(2 downto 0);
signal y_m29b101_1 :  std_logic_vector(2 downto 0);
signal Y0X0_101_m29 :  std_logic_vector(5 downto 0);
signal PP101X0Y0_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w18_0 :  std_logic;
signal heap_bh30_w19_0 :  std_logic;
signal heap_bh30_w20_0 :  std_logic;
signal heap_bh30_w21_0 :  std_logic;
signal heap_bh30_w22_0 :  std_logic;
signal Y0X1_101_m29 :  std_logic_vector(5 downto 0);
signal PP101X1Y0_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w21_1 :  std_logic;
signal heap_bh30_w22_1 :  std_logic;
signal heap_bh30_w23_0 :  std_logic;
signal heap_bh30_w24_0 :  std_logic;
signal heap_bh30_w25_0 :  std_logic;
signal Y0X2_101_m29 :  std_logic_vector(5 downto 0);
signal PP101X2Y0_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w24_1 :  std_logic;
signal heap_bh30_w25_1 :  std_logic;
signal heap_bh30_w26_0 :  std_logic;
signal heap_bh30_w27_0 :  std_logic;
signal heap_bh30_w28_0 :  std_logic;
signal Y0X3_101_m29 :  std_logic_vector(5 downto 0);
signal PP101X3Y0_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w27_1 :  std_logic;
signal heap_bh30_w28_1 :  std_logic;
signal heap_bh30_w29_0 :  std_logic;
signal heap_bh30_w30_0 :  std_logic;
signal heap_bh30_w31_0 :  std_logic;
signal Y0X4_101_m29 :  std_logic_vector(5 downto 0);
signal PP101X4Y0_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w30_1 :  std_logic;
signal heap_bh30_w31_1 :  std_logic;
signal heap_bh30_w32_0 :  std_logic;
signal heap_bh30_w33_0 :  std_logic;
signal heap_bh30_w34_0 :  std_logic;
signal Y0X5_101_m29 :  std_logic_vector(5 downto 0);
signal PP101X5Y0_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w33_1 :  std_logic;
signal heap_bh30_w34_1 :  std_logic;
signal heap_bh30_w35_0 :  std_logic;
signal heap_bh30_w36_0 :  std_logic;
signal heap_bh30_w37_0 :  std_logic;
signal Y0X6_101_m29 :  std_logic_vector(5 downto 0);
signal PP101X6Y0_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w36_1 :  std_logic;
signal heap_bh30_w37_1 :  std_logic;
signal heap_bh30_w38_0 :  std_logic;
signal heap_bh30_w39_0 :  std_logic;
signal heap_bh30_w40_0 :  std_logic;
signal Y0X7_101_m29 :  std_logic_vector(5 downto 0);
signal PP101X7Y0_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w39_1 :  std_logic;
signal heap_bh30_w40_1 :  std_logic;
signal heap_bh30_w41_0 :  std_logic;
signal heap_bh30_w42_1 :  std_logic;
signal heap_bh30_w43_1 :  std_logic;
signal Y1X0_101_m29 :  std_logic_vector(5 downto 0);
signal PP101X0Y1_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w20_1 :  std_logic;
signal heap_bh30_w21_2 :  std_logic;
signal heap_bh30_w22_2 :  std_logic;
signal heap_bh30_w23_1 :  std_logic;
signal heap_bh30_w24_2 :  std_logic;
signal heap_bh30_w25_2 :  std_logic;
signal Y1X1_101_m29 :  std_logic_vector(5 downto 0);
signal PP101X1Y1_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w23_2 :  std_logic;
signal heap_bh30_w24_3 :  std_logic;
signal heap_bh30_w25_3 :  std_logic;
signal heap_bh30_w26_1 :  std_logic;
signal heap_bh30_w27_2 :  std_logic;
signal heap_bh30_w28_2 :  std_logic;
signal Y1X2_101_m29 :  std_logic_vector(5 downto 0);
signal PP101X2Y1_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w26_2 :  std_logic;
signal heap_bh30_w27_3 :  std_logic;
signal heap_bh30_w28_3 :  std_logic;
signal heap_bh30_w29_1 :  std_logic;
signal heap_bh30_w30_2 :  std_logic;
signal heap_bh30_w31_2 :  std_logic;
signal Y1X3_101_m29 :  std_logic_vector(5 downto 0);
signal PP101X3Y1_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w29_2 :  std_logic;
signal heap_bh30_w30_3 :  std_logic;
signal heap_bh30_w31_3 :  std_logic;
signal heap_bh30_w32_1 :  std_logic;
signal heap_bh30_w33_2 :  std_logic;
signal heap_bh30_w34_2 :  std_logic;
signal Y1X4_101_m29 :  std_logic_vector(5 downto 0);
signal PP101X4Y1_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w32_2 :  std_logic;
signal heap_bh30_w33_3 :  std_logic;
signal heap_bh30_w34_3 :  std_logic;
signal heap_bh30_w35_1 :  std_logic;
signal heap_bh30_w36_2 :  std_logic;
signal heap_bh30_w37_2 :  std_logic;
signal Y1X5_101_m29 :  std_logic_vector(5 downto 0);
signal PP101X5Y1_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w35_2 :  std_logic;
signal heap_bh30_w36_3 :  std_logic;
signal heap_bh30_w37_3 :  std_logic;
signal heap_bh30_w38_1 :  std_logic;
signal heap_bh30_w39_2 :  std_logic;
signal heap_bh30_w40_2 :  std_logic;
signal Y1X6_101_m29 :  std_logic_vector(5 downto 0);
signal PP101X6Y1_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w38_2 :  std_logic;
signal heap_bh30_w39_3 :  std_logic;
signal heap_bh30_w40_3 :  std_logic;
signal heap_bh30_w41_1 :  std_logic;
signal heap_bh30_w42_2 :  std_logic;
signal heap_bh30_w43_2 :  std_logic;
signal Y1X7_101_m29 :  std_logic_vector(5 downto 0);
signal PP101X7Y1_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w41_2 :  std_logic;
signal heap_bh30_w42_3 :  std_logic;
signal heap_bh30_w43_3 :  std_logic;
signal heap_bh30_w44_2 :  std_logic;
signal heap_bh30_w45_3 :  std_logic;
signal heap_bh30_w46_3 :  std_logic;
signal Xp_m29b136 :  std_logic_vector(17 downto 0);
signal Yp_m29b136 :  std_logic_vector(5 downto 0);
signal x_m29b136_0 :  std_logic_vector(2 downto 0);
signal x_m29b136_1 :  std_logic_vector(2 downto 0);
signal x_m29b136_2 :  std_logic_vector(2 downto 0);
signal x_m29b136_3 :  std_logic_vector(2 downto 0);
signal x_m29b136_4 :  std_logic_vector(2 downto 0);
signal x_m29b136_5 :  std_logic_vector(2 downto 0);
signal y_m29b136_0 :  std_logic_vector(2 downto 0);
signal y_m29b136_1 :  std_logic_vector(2 downto 0);
signal Y0X0_136_m29 :  std_logic_vector(5 downto 0);
signal PP136X0Y0_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w0_0 :  std_logic;
signal heap_bh30_w1_0 :  std_logic;
signal heap_bh30_w2_0 :  std_logic;
signal heap_bh30_w3_0 :  std_logic;
signal heap_bh30_w4_0 :  std_logic;
signal Y0X1_136_m29 :  std_logic_vector(5 downto 0);
signal PP136X1Y0_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w3_1 :  std_logic;
signal heap_bh30_w4_1 :  std_logic;
signal heap_bh30_w5_0 :  std_logic;
signal heap_bh30_w6_0 :  std_logic;
signal heap_bh30_w7_0 :  std_logic;
signal Y0X2_136_m29 :  std_logic_vector(5 downto 0);
signal PP136X2Y0_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w6_1 :  std_logic;
signal heap_bh30_w7_1 :  std_logic;
signal heap_bh30_w8_0 :  std_logic;
signal heap_bh30_w9_0 :  std_logic;
signal heap_bh30_w10_0 :  std_logic;
signal Y0X3_136_m29 :  std_logic_vector(5 downto 0);
signal PP136X3Y0_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w9_1 :  std_logic;
signal heap_bh30_w10_1 :  std_logic;
signal heap_bh30_w11_0 :  std_logic;
signal heap_bh30_w12_0 :  std_logic;
signal heap_bh30_w13_0 :  std_logic;
signal Y0X4_136_m29 :  std_logic_vector(5 downto 0);
signal PP136X4Y0_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w12_1 :  std_logic;
signal heap_bh30_w13_1 :  std_logic;
signal heap_bh30_w14_0 :  std_logic;
signal heap_bh30_w15_0 :  std_logic;
signal heap_bh30_w16_0 :  std_logic;
signal Y0X5_136_m29 :  std_logic_vector(5 downto 0);
signal PP136X5Y0_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w15_1 :  std_logic;
signal heap_bh30_w16_1 :  std_logic;
signal heap_bh30_w17_0 :  std_logic;
signal heap_bh30_w18_1 :  std_logic;
signal heap_bh30_w19_1 :  std_logic;
signal Y1X0_136_m29 :  std_logic_vector(5 downto 0);
signal PP136X0Y1_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w2_1 :  std_logic;
signal heap_bh30_w3_2 :  std_logic;
signal heap_bh30_w4_2 :  std_logic;
signal heap_bh30_w5_1 :  std_logic;
signal heap_bh30_w6_2 :  std_logic;
signal heap_bh30_w7_2 :  std_logic;
signal Y1X1_136_m29 :  std_logic_vector(5 downto 0);
signal PP136X1Y1_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w5_2 :  std_logic;
signal heap_bh30_w6_3 :  std_logic;
signal heap_bh30_w7_3 :  std_logic;
signal heap_bh30_w8_1 :  std_logic;
signal heap_bh30_w9_2 :  std_logic;
signal heap_bh30_w10_2 :  std_logic;
signal Y1X2_136_m29 :  std_logic_vector(5 downto 0);
signal PP136X2Y1_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w8_2 :  std_logic;
signal heap_bh30_w9_3 :  std_logic;
signal heap_bh30_w10_3 :  std_logic;
signal heap_bh30_w11_1 :  std_logic;
signal heap_bh30_w12_2 :  std_logic;
signal heap_bh30_w13_2 :  std_logic;
signal Y1X3_136_m29 :  std_logic_vector(5 downto 0);
signal PP136X3Y1_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w11_2 :  std_logic;
signal heap_bh30_w12_3 :  std_logic;
signal heap_bh30_w13_3 :  std_logic;
signal heap_bh30_w14_1 :  std_logic;
signal heap_bh30_w15_2 :  std_logic;
signal heap_bh30_w16_2 :  std_logic;
signal Y1X4_136_m29 :  std_logic_vector(5 downto 0);
signal PP136X4Y1_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w14_2 :  std_logic;
signal heap_bh30_w15_3 :  std_logic;
signal heap_bh30_w16_3 :  std_logic;
signal heap_bh30_w17_1 :  std_logic;
signal heap_bh30_w18_2 :  std_logic;
signal heap_bh30_w19_2 :  std_logic;
signal Y1X5_136_m29 :  std_logic_vector(5 downto 0);
signal PP136X5Y1_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w17_2 :  std_logic;
signal heap_bh30_w18_3 :  std_logic;
signal heap_bh30_w19_3 :  std_logic;
signal heap_bh30_w20_2 :  std_logic;
signal heap_bh30_w21_3 :  std_logic;
signal heap_bh30_w22_3 :  std_logic;
signal DSP_bh30_ch0_0 :  std_logic_vector(40 downto 0);
signal heap_bh30_w179_0 :  std_logic;
signal heap_bh30_w178_0 :  std_logic;
signal heap_bh30_w177_0 :  std_logic;
signal heap_bh30_w176_0 :  std_logic;
signal heap_bh30_w175_0 :  std_logic;
signal heap_bh30_w174_0 :  std_logic;
signal heap_bh30_w173_0 :  std_logic;
signal heap_bh30_w172_0 :  std_logic;
signal heap_bh30_w171_0 :  std_logic;
signal heap_bh30_w170_0 :  std_logic;
signal heap_bh30_w169_0 :  std_logic;
signal heap_bh30_w168_0 :  std_logic;
signal heap_bh30_w167_0 :  std_logic;
signal heap_bh30_w166_0 :  std_logic;
signal heap_bh30_w165_0 :  std_logic;
signal heap_bh30_w164_0 :  std_logic;
signal heap_bh30_w163_0 :  std_logic;
signal heap_bh30_w162_0 :  std_logic;
signal heap_bh30_w161_0 :  std_logic;
signal heap_bh30_w160_0 :  std_logic;
signal heap_bh30_w159_0 :  std_logic;
signal heap_bh30_w158_0 :  std_logic;
signal heap_bh30_w157_0 :  std_logic;
signal heap_bh30_w156_0 :  std_logic;
signal heap_bh30_w155_0 :  std_logic;
signal heap_bh30_w154_0 :  std_logic;
signal heap_bh30_w153_0 :  std_logic;
signal heap_bh30_w152_0 :  std_logic;
signal heap_bh30_w151_0 :  std_logic;
signal heap_bh30_w150_0 :  std_logic;
signal heap_bh30_w149_0 :  std_logic;
signal heap_bh30_w148_0 :  std_logic;
signal heap_bh30_w147_0 :  std_logic;
signal heap_bh30_w146_0 :  std_logic;
signal heap_bh30_w145_0 :  std_logic;
signal heap_bh30_w144_0 :  std_logic;
signal heap_bh30_w143_0 :  std_logic;
signal heap_bh30_w142_0 :  std_logic;
signal heap_bh30_w141_0 :  std_logic;
signal heap_bh30_w140_0 :  std_logic;
signal heap_bh30_w139_0 :  std_logic;
signal DSP_bh30_ch1_0 :  std_logic_vector(40 downto 0);
signal heap_bh30_w155_1 :  std_logic;
signal heap_bh30_w154_1 :  std_logic;
signal heap_bh30_w153_1 :  std_logic;
signal heap_bh30_w152_1 :  std_logic;
signal heap_bh30_w151_1 :  std_logic;
signal heap_bh30_w150_1 :  std_logic;
signal heap_bh30_w149_1 :  std_logic;
signal heap_bh30_w148_1 :  std_logic;
signal heap_bh30_w147_1 :  std_logic;
signal heap_bh30_w146_1 :  std_logic;
signal heap_bh30_w145_1 :  std_logic;
signal heap_bh30_w144_1 :  std_logic;
signal heap_bh30_w143_1 :  std_logic;
signal heap_bh30_w142_1 :  std_logic;
signal heap_bh30_w141_1 :  std_logic;
signal heap_bh30_w140_1 :  std_logic;
signal heap_bh30_w139_1 :  std_logic;
signal heap_bh30_w138_0 :  std_logic;
signal heap_bh30_w137_0 :  std_logic;
signal heap_bh30_w136_0 :  std_logic;
signal heap_bh30_w135_0 :  std_logic;
signal heap_bh30_w134_0 :  std_logic;
signal heap_bh30_w133_0 :  std_logic;
signal heap_bh30_w132_0 :  std_logic;
signal heap_bh30_w131_0 :  std_logic;
signal heap_bh30_w130_0 :  std_logic;
signal heap_bh30_w129_0 :  std_logic;
signal heap_bh30_w128_0 :  std_logic;
signal heap_bh30_w127_0 :  std_logic;
signal heap_bh30_w126_0 :  std_logic;
signal heap_bh30_w125_0 :  std_logic;
signal heap_bh30_w124_0 :  std_logic;
signal heap_bh30_w123_0 :  std_logic;
signal heap_bh30_w122_0 :  std_logic;
signal heap_bh30_w121_0 :  std_logic;
signal heap_bh30_w120_0 :  std_logic;
signal heap_bh30_w119_0 :  std_logic;
signal heap_bh30_w118_0 :  std_logic;
signal heap_bh30_w117_0 :  std_logic;
signal heap_bh30_w116_0 :  std_logic;
signal heap_bh30_w115_0 :  std_logic;
signal DSP_bh30_ch2_0 :  std_logic_vector(40 downto 0);
signal heap_bh30_w131_1 :  std_logic;
signal heap_bh30_w130_1 :  std_logic;
signal heap_bh30_w129_1 :  std_logic;
signal heap_bh30_w128_1 :  std_logic;
signal heap_bh30_w127_1 :  std_logic;
signal heap_bh30_w126_1 :  std_logic;
signal heap_bh30_w125_1 :  std_logic;
signal heap_bh30_w124_1 :  std_logic;
signal heap_bh30_w123_1 :  std_logic;
signal heap_bh30_w122_1 :  std_logic;
signal heap_bh30_w121_1 :  std_logic;
signal heap_bh30_w120_1 :  std_logic;
signal heap_bh30_w119_1 :  std_logic;
signal heap_bh30_w118_1 :  std_logic;
signal heap_bh30_w117_1 :  std_logic;
signal heap_bh30_w116_1 :  std_logic;
signal heap_bh30_w115_1 :  std_logic;
signal heap_bh30_w114_0 :  std_logic;
signal heap_bh30_w113_0 :  std_logic;
signal heap_bh30_w112_0 :  std_logic;
signal heap_bh30_w111_0 :  std_logic;
signal heap_bh30_w110_0 :  std_logic;
signal heap_bh30_w109_0 :  std_logic;
signal heap_bh30_w108_0 :  std_logic;
signal heap_bh30_w107_0 :  std_logic;
signal heap_bh30_w106_0 :  std_logic;
signal heap_bh30_w105_0 :  std_logic;
signal heap_bh30_w104_0 :  std_logic;
signal heap_bh30_w103_0 :  std_logic;
signal heap_bh30_w102_0 :  std_logic;
signal heap_bh30_w101_0 :  std_logic;
signal heap_bh30_w100_0 :  std_logic;
signal heap_bh30_w99_0 :  std_logic;
signal heap_bh30_w98_0 :  std_logic;
signal heap_bh30_w97_0 :  std_logic;
signal heap_bh30_w96_0 :  std_logic;
signal heap_bh30_w95_0 :  std_logic;
signal heap_bh30_w94_1 :  std_logic;
signal heap_bh30_w93_1 :  std_logic;
signal heap_bh30_w92_1 :  std_logic;
signal heap_bh30_w91_3 :  std_logic;
signal DSP_bh30_ch3_0 :  std_logic_vector(40 downto 0);
signal heap_bh30_w107_1 :  std_logic;
signal heap_bh30_w106_1 :  std_logic;
signal heap_bh30_w105_1 :  std_logic;
signal heap_bh30_w104_1 :  std_logic;
signal heap_bh30_w103_1 :  std_logic;
signal heap_bh30_w102_1 :  std_logic;
signal heap_bh30_w101_1 :  std_logic;
signal heap_bh30_w100_1 :  std_logic;
signal heap_bh30_w99_1 :  std_logic;
signal heap_bh30_w98_1 :  std_logic;
signal heap_bh30_w97_1 :  std_logic;
signal heap_bh30_w96_1 :  std_logic;
signal heap_bh30_w95_1 :  std_logic;
signal heap_bh30_w94_2 :  std_logic;
signal heap_bh30_w93_2 :  std_logic;
signal heap_bh30_w92_2 :  std_logic;
signal heap_bh30_w91_4 :  std_logic;
signal heap_bh30_w90_3 :  std_logic;
signal heap_bh30_w89_3 :  std_logic;
signal heap_bh30_w88_4 :  std_logic;
signal heap_bh30_w87_4 :  std_logic;
signal heap_bh30_w86_3 :  std_logic;
signal heap_bh30_w85_4 :  std_logic;
signal heap_bh30_w84_4 :  std_logic;
signal heap_bh30_w83_3 :  std_logic;
signal heap_bh30_w82_4 :  std_logic;
signal heap_bh30_w81_4 :  std_logic;
signal heap_bh30_w80_3 :  std_logic;
signal heap_bh30_w79_4 :  std_logic;
signal heap_bh30_w78_4 :  std_logic;
signal heap_bh30_w77_3 :  std_logic;
signal heap_bh30_w76_4 :  std_logic;
signal heap_bh30_w75_4 :  std_logic;
signal heap_bh30_w74_3 :  std_logic;
signal heap_bh30_w73_4 :  std_logic;
signal heap_bh30_w72_4 :  std_logic;
signal heap_bh30_w71_3 :  std_logic;
signal heap_bh30_w70_4 :  std_logic;
signal heap_bh30_w69_4 :  std_logic;
signal heap_bh30_w68_3 :  std_logic;
signal heap_bh30_w67_4 :  std_logic;
signal DSP_bh30_ch4_0 :  std_logic_vector(40 downto 0);
signal heap_bh30_w162_1 :  std_logic;
signal heap_bh30_w161_1 :  std_logic;
signal heap_bh30_w160_1 :  std_logic;
signal heap_bh30_w159_1 :  std_logic;
signal heap_bh30_w158_1 :  std_logic;
signal heap_bh30_w157_1 :  std_logic;
signal heap_bh30_w156_1 :  std_logic;
signal heap_bh30_w155_2 :  std_logic;
signal heap_bh30_w154_2 :  std_logic;
signal heap_bh30_w153_2 :  std_logic;
signal heap_bh30_w152_2 :  std_logic;
signal heap_bh30_w151_2 :  std_logic;
signal heap_bh30_w150_2 :  std_logic;
signal heap_bh30_w149_2 :  std_logic;
signal heap_bh30_w148_2 :  std_logic;
signal heap_bh30_w147_2 :  std_logic;
signal heap_bh30_w146_2 :  std_logic;
signal heap_bh30_w145_2 :  std_logic;
signal heap_bh30_w144_2 :  std_logic;
signal heap_bh30_w143_2 :  std_logic;
signal heap_bh30_w142_2 :  std_logic;
signal heap_bh30_w141_2 :  std_logic;
signal heap_bh30_w140_2 :  std_logic;
signal heap_bh30_w139_2 :  std_logic;
signal heap_bh30_w138_1 :  std_logic;
signal heap_bh30_w137_1 :  std_logic;
signal heap_bh30_w136_1 :  std_logic;
signal heap_bh30_w135_1 :  std_logic;
signal heap_bh30_w134_1 :  std_logic;
signal heap_bh30_w133_1 :  std_logic;
signal heap_bh30_w132_1 :  std_logic;
signal heap_bh30_w131_2 :  std_logic;
signal heap_bh30_w130_2 :  std_logic;
signal heap_bh30_w129_2 :  std_logic;
signal heap_bh30_w128_2 :  std_logic;
signal heap_bh30_w127_2 :  std_logic;
signal heap_bh30_w126_2 :  std_logic;
signal heap_bh30_w125_2 :  std_logic;
signal heap_bh30_w124_2 :  std_logic;
signal heap_bh30_w123_2 :  std_logic;
signal heap_bh30_w122_2 :  std_logic;
signal DSP_bh30_ch5_0 :  std_logic_vector(40 downto 0);
signal heap_bh30_w138_2 :  std_logic;
signal heap_bh30_w137_2 :  std_logic;
signal heap_bh30_w136_2 :  std_logic;
signal heap_bh30_w135_2 :  std_logic;
signal heap_bh30_w134_2 :  std_logic;
signal heap_bh30_w133_2 :  std_logic;
signal heap_bh30_w132_2 :  std_logic;
signal heap_bh30_w131_3 :  std_logic;
signal heap_bh30_w130_3 :  std_logic;
signal heap_bh30_w129_3 :  std_logic;
signal heap_bh30_w128_3 :  std_logic;
signal heap_bh30_w127_3 :  std_logic;
signal heap_bh30_w126_3 :  std_logic;
signal heap_bh30_w125_3 :  std_logic;
signal heap_bh30_w124_3 :  std_logic;
signal heap_bh30_w123_3 :  std_logic;
signal heap_bh30_w122_3 :  std_logic;
signal heap_bh30_w121_2 :  std_logic;
signal heap_bh30_w120_2 :  std_logic;
signal heap_bh30_w119_2 :  std_logic;
signal heap_bh30_w118_2 :  std_logic;
signal heap_bh30_w117_2 :  std_logic;
signal heap_bh30_w116_2 :  std_logic;
signal heap_bh30_w115_2 :  std_logic;
signal heap_bh30_w114_1 :  std_logic;
signal heap_bh30_w113_1 :  std_logic;
signal heap_bh30_w112_1 :  std_logic;
signal heap_bh30_w111_1 :  std_logic;
signal heap_bh30_w110_1 :  std_logic;
signal heap_bh30_w109_1 :  std_logic;
signal heap_bh30_w108_1 :  std_logic;
signal heap_bh30_w107_2 :  std_logic;
signal heap_bh30_w106_2 :  std_logic;
signal heap_bh30_w105_2 :  std_logic;
signal heap_bh30_w104_2 :  std_logic;
signal heap_bh30_w103_2 :  std_logic;
signal heap_bh30_w102_2 :  std_logic;
signal heap_bh30_w101_2 :  std_logic;
signal heap_bh30_w100_2 :  std_logic;
signal heap_bh30_w99_2 :  std_logic;
signal heap_bh30_w98_2 :  std_logic;
signal DSP_bh30_ch6_0 :  std_logic_vector(40 downto 0);
signal heap_bh30_w114_2 :  std_logic;
signal heap_bh30_w113_2 :  std_logic;
signal heap_bh30_w112_2 :  std_logic;
signal heap_bh30_w111_2 :  std_logic;
signal heap_bh30_w110_2 :  std_logic;
signal heap_bh30_w109_2 :  std_logic;
signal heap_bh30_w108_2 :  std_logic;
signal heap_bh30_w107_3 :  std_logic;
signal heap_bh30_w106_3 :  std_logic;
signal heap_bh30_w105_3 :  std_logic;
signal heap_bh30_w104_3 :  std_logic;
signal heap_bh30_w103_3 :  std_logic;
signal heap_bh30_w102_3 :  std_logic;
signal heap_bh30_w101_3 :  std_logic;
signal heap_bh30_w100_3 :  std_logic;
signal heap_bh30_w99_3 :  std_logic;
signal heap_bh30_w98_3 :  std_logic;
signal heap_bh30_w97_2 :  std_logic;
signal heap_bh30_w96_2 :  std_logic;
signal heap_bh30_w95_2 :  std_logic;
signal heap_bh30_w94_3 :  std_logic;
signal heap_bh30_w93_3 :  std_logic;
signal heap_bh30_w92_3 :  std_logic;
signal heap_bh30_w91_5 :  std_logic;
signal heap_bh30_w90_4 :  std_logic;
signal heap_bh30_w89_4 :  std_logic;
signal heap_bh30_w88_5 :  std_logic;
signal heap_bh30_w87_5 :  std_logic;
signal heap_bh30_w86_4 :  std_logic;
signal heap_bh30_w85_5 :  std_logic;
signal heap_bh30_w84_5 :  std_logic;
signal heap_bh30_w83_4 :  std_logic;
signal heap_bh30_w82_5 :  std_logic;
signal heap_bh30_w81_5 :  std_logic;
signal heap_bh30_w80_4 :  std_logic;
signal heap_bh30_w79_5 :  std_logic;
signal heap_bh30_w78_5 :  std_logic;
signal heap_bh30_w77_4 :  std_logic;
signal heap_bh30_w76_5 :  std_logic;
signal heap_bh30_w75_5 :  std_logic;
signal heap_bh30_w74_4 :  std_logic;
signal DSP_bh30_ch7_0 :  std_logic_vector(40 downto 0);
signal heap_bh30_w90_5 :  std_logic;
signal heap_bh30_w89_5 :  std_logic;
signal heap_bh30_w88_6 :  std_logic;
signal heap_bh30_w87_6 :  std_logic;
signal heap_bh30_w86_5 :  std_logic;
signal heap_bh30_w85_6 :  std_logic;
signal heap_bh30_w84_6 :  std_logic;
signal heap_bh30_w83_5 :  std_logic;
signal heap_bh30_w82_6 :  std_logic;
signal heap_bh30_w81_6 :  std_logic;
signal heap_bh30_w80_5 :  std_logic;
signal heap_bh30_w79_6 :  std_logic;
signal heap_bh30_w78_6 :  std_logic;
signal heap_bh30_w77_5 :  std_logic;
signal heap_bh30_w76_6 :  std_logic;
signal heap_bh30_w75_6 :  std_logic;
signal heap_bh30_w74_5 :  std_logic;
signal heap_bh30_w73_5 :  std_logic;
signal heap_bh30_w72_5 :  std_logic;
signal heap_bh30_w71_4 :  std_logic;
signal heap_bh30_w70_5 :  std_logic;
signal heap_bh30_w69_5 :  std_logic;
signal heap_bh30_w68_4 :  std_logic;
signal heap_bh30_w67_5 :  std_logic;
signal heap_bh30_w66_4 :  std_logic;
signal heap_bh30_w65_3 :  std_logic;
signal heap_bh30_w64_4 :  std_logic;
signal heap_bh30_w63_4 :  std_logic;
signal heap_bh30_w62_3 :  std_logic;
signal heap_bh30_w61_4 :  std_logic;
signal heap_bh30_w60_4 :  std_logic;
signal heap_bh30_w59_3 :  std_logic;
signal heap_bh30_w58_4 :  std_logic;
signal heap_bh30_w57_4 :  std_logic;
signal heap_bh30_w56_3 :  std_logic;
signal heap_bh30_w55_4 :  std_logic;
signal heap_bh30_w54_4 :  std_logic;
signal heap_bh30_w53_3 :  std_logic;
signal heap_bh30_w52_4 :  std_logic;
signal heap_bh30_w51_4 :  std_logic;
signal heap_bh30_w50_3 :  std_logic;
signal DSP_bh30_ch8_0 :  std_logic_vector(40 downto 0);
signal heap_bh30_w145_3 :  std_logic;
signal heap_bh30_w144_3 :  std_logic;
signal heap_bh30_w143_3 :  std_logic;
signal heap_bh30_w142_3 :  std_logic;
signal heap_bh30_w141_3 :  std_logic;
signal heap_bh30_w140_3 :  std_logic;
signal heap_bh30_w139_3 :  std_logic;
signal heap_bh30_w138_3 :  std_logic;
signal heap_bh30_w137_3 :  std_logic;
signal heap_bh30_w136_3 :  std_logic;
signal heap_bh30_w135_3 :  std_logic;
signal heap_bh30_w134_3 :  std_logic;
signal heap_bh30_w133_3 :  std_logic;
signal heap_bh30_w132_3 :  std_logic;
signal heap_bh30_w131_4 :  std_logic;
signal heap_bh30_w130_4 :  std_logic;
signal heap_bh30_w129_4 :  std_logic;
signal heap_bh30_w128_4 :  std_logic;
signal heap_bh30_w127_4 :  std_logic;
signal heap_bh30_w126_4 :  std_logic;
signal heap_bh30_w125_4 :  std_logic;
signal heap_bh30_w124_4 :  std_logic;
signal heap_bh30_w123_4 :  std_logic;
signal heap_bh30_w122_4 :  std_logic;
signal heap_bh30_w121_3 :  std_logic;
signal heap_bh30_w120_3 :  std_logic;
signal heap_bh30_w119_3 :  std_logic;
signal heap_bh30_w118_3 :  std_logic;
signal heap_bh30_w117_3 :  std_logic;
signal heap_bh30_w116_3 :  std_logic;
signal heap_bh30_w115_3 :  std_logic;
signal heap_bh30_w114_3 :  std_logic;
signal heap_bh30_w113_3 :  std_logic;
signal heap_bh30_w112_3 :  std_logic;
signal heap_bh30_w111_3 :  std_logic;
signal heap_bh30_w110_3 :  std_logic;
signal heap_bh30_w109_3 :  std_logic;
signal heap_bh30_w108_3 :  std_logic;
signal heap_bh30_w107_4 :  std_logic;
signal heap_bh30_w106_4 :  std_logic;
signal heap_bh30_w105_4 :  std_logic;
signal DSP_bh30_ch9_0 :  std_logic_vector(40 downto 0);
signal heap_bh30_w121_4 :  std_logic;
signal heap_bh30_w120_4 :  std_logic;
signal heap_bh30_w119_4 :  std_logic;
signal heap_bh30_w118_4 :  std_logic;
signal heap_bh30_w117_4 :  std_logic;
signal heap_bh30_w116_4 :  std_logic;
signal heap_bh30_w115_4 :  std_logic;
signal heap_bh30_w114_4 :  std_logic;
signal heap_bh30_w113_4 :  std_logic;
signal heap_bh30_w112_4 :  std_logic;
signal heap_bh30_w111_4 :  std_logic;
signal heap_bh30_w110_4 :  std_logic;
signal heap_bh30_w109_4 :  std_logic;
signal heap_bh30_w108_4 :  std_logic;
signal heap_bh30_w107_5 :  std_logic;
signal heap_bh30_w106_5 :  std_logic;
signal heap_bh30_w105_5 :  std_logic;
signal heap_bh30_w104_4 :  std_logic;
signal heap_bh30_w103_4 :  std_logic;
signal heap_bh30_w102_4 :  std_logic;
signal heap_bh30_w101_4 :  std_logic;
signal heap_bh30_w100_4 :  std_logic;
signal heap_bh30_w99_4 :  std_logic;
signal heap_bh30_w98_4 :  std_logic;
signal heap_bh30_w97_3 :  std_logic;
signal heap_bh30_w96_3 :  std_logic;
signal heap_bh30_w95_3 :  std_logic;
signal heap_bh30_w94_4 :  std_logic;
signal heap_bh30_w93_4 :  std_logic;
signal heap_bh30_w92_4 :  std_logic;
signal heap_bh30_w91_6 :  std_logic;
signal heap_bh30_w90_6 :  std_logic;
signal heap_bh30_w89_6 :  std_logic;
signal heap_bh30_w88_7 :  std_logic;
signal heap_bh30_w87_7 :  std_logic;
signal heap_bh30_w86_6 :  std_logic;
signal heap_bh30_w85_7 :  std_logic;
signal heap_bh30_w84_7 :  std_logic;
signal heap_bh30_w83_6 :  std_logic;
signal heap_bh30_w82_7 :  std_logic;
signal heap_bh30_w81_7 :  std_logic;
signal DSP_bh30_ch10_0 :  std_logic_vector(40 downto 0);
signal heap_bh30_w97_4 :  std_logic;
signal heap_bh30_w96_4 :  std_logic;
signal heap_bh30_w95_4 :  std_logic;
signal heap_bh30_w94_5 :  std_logic;
signal heap_bh30_w93_5 :  std_logic;
signal heap_bh30_w92_5 :  std_logic;
signal heap_bh30_w91_7 :  std_logic;
signal heap_bh30_w90_7 :  std_logic;
signal heap_bh30_w89_7 :  std_logic;
signal heap_bh30_w88_8 :  std_logic;
signal heap_bh30_w87_8 :  std_logic;
signal heap_bh30_w86_7 :  std_logic;
signal heap_bh30_w85_8 :  std_logic;
signal heap_bh30_w84_8 :  std_logic;
signal heap_bh30_w83_7 :  std_logic;
signal heap_bh30_w82_8 :  std_logic;
signal heap_bh30_w81_8 :  std_logic;
signal heap_bh30_w80_6 :  std_logic;
signal heap_bh30_w79_7 :  std_logic;
signal heap_bh30_w78_7 :  std_logic;
signal heap_bh30_w77_6 :  std_logic;
signal heap_bh30_w76_7 :  std_logic;
signal heap_bh30_w75_7 :  std_logic;
signal heap_bh30_w74_6 :  std_logic;
signal heap_bh30_w73_6 :  std_logic;
signal heap_bh30_w72_6 :  std_logic;
signal heap_bh30_w71_5 :  std_logic;
signal heap_bh30_w70_6 :  std_logic;
signal heap_bh30_w69_6 :  std_logic;
signal heap_bh30_w68_5 :  std_logic;
signal heap_bh30_w67_6 :  std_logic;
signal heap_bh30_w66_5 :  std_logic;
signal heap_bh30_w65_4 :  std_logic;
signal heap_bh30_w64_5 :  std_logic;
signal heap_bh30_w63_5 :  std_logic;
signal heap_bh30_w62_4 :  std_logic;
signal heap_bh30_w61_5 :  std_logic;
signal heap_bh30_w60_5 :  std_logic;
signal heap_bh30_w59_4 :  std_logic;
signal heap_bh30_w58_5 :  std_logic;
signal heap_bh30_w57_5 :  std_logic;
signal DSP_bh30_ch11_0 :  std_logic_vector(40 downto 0);
signal heap_bh30_w73_7 :  std_logic;
signal heap_bh30_w72_7 :  std_logic;
signal heap_bh30_w71_6 :  std_logic;
signal heap_bh30_w70_7 :  std_logic;
signal heap_bh30_w69_7 :  std_logic;
signal heap_bh30_w68_6 :  std_logic;
signal heap_bh30_w67_7 :  std_logic;
signal heap_bh30_w66_6 :  std_logic;
signal heap_bh30_w65_5 :  std_logic;
signal heap_bh30_w64_6 :  std_logic;
signal heap_bh30_w63_6 :  std_logic;
signal heap_bh30_w62_5 :  std_logic;
signal heap_bh30_w61_6 :  std_logic;
signal heap_bh30_w60_6 :  std_logic;
signal heap_bh30_w59_5 :  std_logic;
signal heap_bh30_w58_6 :  std_logic;
signal heap_bh30_w57_6 :  std_logic;
signal heap_bh30_w56_4 :  std_logic;
signal heap_bh30_w55_5 :  std_logic;
signal heap_bh30_w54_5 :  std_logic;
signal heap_bh30_w53_4 :  std_logic;
signal heap_bh30_w52_5 :  std_logic;
signal heap_bh30_w51_5 :  std_logic;
signal heap_bh30_w50_4 :  std_logic;
signal heap_bh30_w49_4 :  std_logic;
signal heap_bh30_w48_4 :  std_logic;
signal heap_bh30_w47_3 :  std_logic;
signal heap_bh30_w46_4 :  std_logic;
signal heap_bh30_w45_4 :  std_logic;
signal heap_bh30_w44_3 :  std_logic;
signal heap_bh30_w43_4 :  std_logic;
signal heap_bh30_w42_4 :  std_logic;
signal heap_bh30_w41_3 :  std_logic;
signal heap_bh30_w40_4 :  std_logic;
signal heap_bh30_w39_4 :  std_logic;
signal heap_bh30_w38_3 :  std_logic;
signal heap_bh30_w37_4 :  std_logic;
signal heap_bh30_w36_4 :  std_logic;
signal heap_bh30_w35_3 :  std_logic;
signal heap_bh30_w34_4 :  std_logic;
signal heap_bh30_w33_4 :  std_logic;
signal DSP_bh30_ch12_0 :  std_logic_vector(40 downto 0);
signal heap_bh30_w128_5 :  std_logic;
signal heap_bh30_w127_5 :  std_logic;
signal heap_bh30_w126_5 :  std_logic;
signal heap_bh30_w125_5 :  std_logic;
signal heap_bh30_w124_5 :  std_logic;
signal heap_bh30_w123_5 :  std_logic;
signal heap_bh30_w122_5 :  std_logic;
signal heap_bh30_w121_5 :  std_logic;
signal heap_bh30_w120_5 :  std_logic;
signal heap_bh30_w119_5 :  std_logic;
signal heap_bh30_w118_5 :  std_logic;
signal heap_bh30_w117_5 :  std_logic;
signal heap_bh30_w116_5 :  std_logic;
signal heap_bh30_w115_5 :  std_logic;
signal heap_bh30_w114_5 :  std_logic;
signal heap_bh30_w113_5 :  std_logic;
signal heap_bh30_w112_5 :  std_logic;
signal heap_bh30_w111_5 :  std_logic;
signal heap_bh30_w110_5 :  std_logic;
signal heap_bh30_w109_5 :  std_logic;
signal heap_bh30_w108_5 :  std_logic;
signal heap_bh30_w107_6 :  std_logic;
signal heap_bh30_w106_6 :  std_logic;
signal heap_bh30_w105_6 :  std_logic;
signal heap_bh30_w104_5 :  std_logic;
signal heap_bh30_w103_5 :  std_logic;
signal heap_bh30_w102_5 :  std_logic;
signal heap_bh30_w101_5 :  std_logic;
signal heap_bh30_w100_5 :  std_logic;
signal heap_bh30_w99_5 :  std_logic;
signal heap_bh30_w98_5 :  std_logic;
signal heap_bh30_w97_5 :  std_logic;
signal heap_bh30_w96_5 :  std_logic;
signal heap_bh30_w95_5 :  std_logic;
signal heap_bh30_w94_6 :  std_logic;
signal heap_bh30_w93_6 :  std_logic;
signal heap_bh30_w92_6 :  std_logic;
signal heap_bh30_w91_8 :  std_logic;
signal heap_bh30_w90_8 :  std_logic;
signal heap_bh30_w89_8 :  std_logic;
signal heap_bh30_w88_9 :  std_logic;
signal DSP_bh30_ch13_0 :  std_logic_vector(40 downto 0);
signal heap_bh30_w104_6 :  std_logic;
signal heap_bh30_w103_6 :  std_logic;
signal heap_bh30_w102_6 :  std_logic;
signal heap_bh30_w101_6 :  std_logic;
signal heap_bh30_w100_6 :  std_logic;
signal heap_bh30_w99_6 :  std_logic;
signal heap_bh30_w98_6 :  std_logic;
signal heap_bh30_w97_6 :  std_logic;
signal heap_bh30_w96_6 :  std_logic;
signal heap_bh30_w95_6 :  std_logic;
signal heap_bh30_w94_7 :  std_logic;
signal heap_bh30_w93_7 :  std_logic;
signal heap_bh30_w92_7 :  std_logic;
signal heap_bh30_w91_9 :  std_logic;
signal heap_bh30_w90_9 :  std_logic;
signal heap_bh30_w89_9 :  std_logic;
signal heap_bh30_w88_10 :  std_logic;
signal heap_bh30_w87_9 :  std_logic;
signal heap_bh30_w86_8 :  std_logic;
signal heap_bh30_w85_9 :  std_logic;
signal heap_bh30_w84_9 :  std_logic;
signal heap_bh30_w83_8 :  std_logic;
signal heap_bh30_w82_9 :  std_logic;
signal heap_bh30_w81_9 :  std_logic;
signal heap_bh30_w80_7 :  std_logic;
signal heap_bh30_w79_8 :  std_logic;
signal heap_bh30_w78_8 :  std_logic;
signal heap_bh30_w77_7 :  std_logic;
signal heap_bh30_w76_8 :  std_logic;
signal heap_bh30_w75_8 :  std_logic;
signal heap_bh30_w74_7 :  std_logic;
signal heap_bh30_w73_8 :  std_logic;
signal heap_bh30_w72_8 :  std_logic;
signal heap_bh30_w71_7 :  std_logic;
signal heap_bh30_w70_8 :  std_logic;
signal heap_bh30_w69_8 :  std_logic;
signal heap_bh30_w68_7 :  std_logic;
signal heap_bh30_w67_8 :  std_logic;
signal heap_bh30_w66_7 :  std_logic;
signal heap_bh30_w65_6 :  std_logic;
signal heap_bh30_w64_7 :  std_logic;
signal DSP_bh30_ch14_0 :  std_logic_vector(40 downto 0);
signal heap_bh30_w80_8 :  std_logic;
signal heap_bh30_w79_9 :  std_logic;
signal heap_bh30_w78_9 :  std_logic;
signal heap_bh30_w77_8 :  std_logic;
signal heap_bh30_w76_9 :  std_logic;
signal heap_bh30_w75_9 :  std_logic;
signal heap_bh30_w74_8 :  std_logic;
signal heap_bh30_w73_9 :  std_logic;
signal heap_bh30_w72_9 :  std_logic;
signal heap_bh30_w71_8 :  std_logic;
signal heap_bh30_w70_9 :  std_logic;
signal heap_bh30_w69_9 :  std_logic;
signal heap_bh30_w68_8 :  std_logic;
signal heap_bh30_w67_9 :  std_logic;
signal heap_bh30_w66_8 :  std_logic;
signal heap_bh30_w65_7 :  std_logic;
signal heap_bh30_w64_8 :  std_logic;
signal heap_bh30_w63_7 :  std_logic;
signal heap_bh30_w62_6 :  std_logic;
signal heap_bh30_w61_7 :  std_logic;
signal heap_bh30_w60_7 :  std_logic;
signal heap_bh30_w59_6 :  std_logic;
signal heap_bh30_w58_7 :  std_logic;
signal heap_bh30_w57_7 :  std_logic;
signal heap_bh30_w56_5 :  std_logic;
signal heap_bh30_w55_6 :  std_logic;
signal heap_bh30_w54_6 :  std_logic;
signal heap_bh30_w53_5 :  std_logic;
signal heap_bh30_w52_6 :  std_logic;
signal heap_bh30_w51_6 :  std_logic;
signal heap_bh30_w50_5 :  std_logic;
signal heap_bh30_w49_5 :  std_logic;
signal heap_bh30_w48_5 :  std_logic;
signal heap_bh30_w47_4 :  std_logic;
signal heap_bh30_w46_5 :  std_logic;
signal heap_bh30_w45_5 :  std_logic;
signal heap_bh30_w44_4 :  std_logic;
signal heap_bh30_w43_5 :  std_logic;
signal heap_bh30_w42_5 :  std_logic;
signal heap_bh30_w41_4 :  std_logic;
signal heap_bh30_w40_5 :  std_logic;
signal DSP_bh30_ch15_0 :  std_logic_vector(40 downto 0);
signal heap_bh30_w56_6 :  std_logic;
signal heap_bh30_w55_7 :  std_logic;
signal heap_bh30_w54_7 :  std_logic;
signal heap_bh30_w53_6 :  std_logic;
signal heap_bh30_w52_7 :  std_logic;
signal heap_bh30_w51_7 :  std_logic;
signal heap_bh30_w50_6 :  std_logic;
signal heap_bh30_w49_6 :  std_logic;
signal heap_bh30_w48_6 :  std_logic;
signal heap_bh30_w47_5 :  std_logic;
signal heap_bh30_w46_6 :  std_logic;
signal heap_bh30_w45_6 :  std_logic;
signal heap_bh30_w44_5 :  std_logic;
signal heap_bh30_w43_6 :  std_logic;
signal heap_bh30_w42_6 :  std_logic;
signal heap_bh30_w41_5 :  std_logic;
signal heap_bh30_w40_6 :  std_logic;
signal heap_bh30_w39_5 :  std_logic;
signal heap_bh30_w38_4 :  std_logic;
signal heap_bh30_w37_5 :  std_logic;
signal heap_bh30_w36_5 :  std_logic;
signal heap_bh30_w35_4 :  std_logic;
signal heap_bh30_w34_5 :  std_logic;
signal heap_bh30_w33_5 :  std_logic;
signal heap_bh30_w32_3 :  std_logic;
signal heap_bh30_w31_4 :  std_logic;
signal heap_bh30_w30_4 :  std_logic;
signal heap_bh30_w29_3 :  std_logic;
signal heap_bh30_w28_4 :  std_logic;
signal heap_bh30_w27_4 :  std_logic;
signal heap_bh30_w26_3 :  std_logic;
signal heap_bh30_w25_4 :  std_logic;
signal heap_bh30_w24_4 :  std_logic;
signal heap_bh30_w23_3 :  std_logic;
signal heap_bh30_w22_4 :  std_logic;
signal heap_bh30_w21_4 :  std_logic;
signal heap_bh30_w20_3 :  std_logic;
signal heap_bh30_w19_4 :  std_logic;
signal heap_bh30_w18_4 :  std_logic;
signal heap_bh30_w17_3 :  std_logic;
signal heap_bh30_w16_4 :  std_logic;
signal DSP_bh30_ch16_0 :  std_logic_vector(40 downto 0);
signal heap_bh30_w111_6 :  std_logic;
signal heap_bh30_w110_6 :  std_logic;
signal heap_bh30_w109_6 :  std_logic;
signal heap_bh30_w108_6 :  std_logic;
signal heap_bh30_w107_7 :  std_logic;
signal heap_bh30_w106_7 :  std_logic;
signal heap_bh30_w105_7 :  std_logic;
signal heap_bh30_w104_7 :  std_logic;
signal heap_bh30_w103_7 :  std_logic;
signal heap_bh30_w102_7 :  std_logic;
signal heap_bh30_w101_7 :  std_logic;
signal heap_bh30_w100_7 :  std_logic;
signal heap_bh30_w99_7 :  std_logic;
signal heap_bh30_w98_7 :  std_logic;
signal heap_bh30_w97_7 :  std_logic;
signal heap_bh30_w96_7 :  std_logic;
signal heap_bh30_w95_7 :  std_logic;
signal heap_bh30_w94_8 :  std_logic;
signal heap_bh30_w93_8 :  std_logic;
signal heap_bh30_w92_8 :  std_logic;
signal heap_bh30_w91_10 :  std_logic;
signal heap_bh30_w90_10 :  std_logic;
signal heap_bh30_w89_10 :  std_logic;
signal heap_bh30_w88_11 :  std_logic;
signal heap_bh30_w87_10 :  std_logic;
signal heap_bh30_w86_9 :  std_logic;
signal heap_bh30_w85_10 :  std_logic;
signal heap_bh30_w84_10 :  std_logic;
signal heap_bh30_w83_9 :  std_logic;
signal heap_bh30_w82_10 :  std_logic;
signal heap_bh30_w81_10 :  std_logic;
signal heap_bh30_w80_9 :  std_logic;
signal heap_bh30_w79_10 :  std_logic;
signal heap_bh30_w78_10 :  std_logic;
signal heap_bh30_w77_9 :  std_logic;
signal heap_bh30_w76_10 :  std_logic;
signal heap_bh30_w75_10 :  std_logic;
signal heap_bh30_w74_9 :  std_logic;
signal heap_bh30_w73_10 :  std_logic;
signal heap_bh30_w72_10 :  std_logic;
signal heap_bh30_w71_9 :  std_logic;
signal DSP_bh30_ch17_0 :  std_logic_vector(40 downto 0);
signal heap_bh30_w87_11 :  std_logic;
signal heap_bh30_w86_10 :  std_logic;
signal heap_bh30_w85_11 :  std_logic;
signal heap_bh30_w84_11 :  std_logic;
signal heap_bh30_w83_10 :  std_logic;
signal heap_bh30_w82_11 :  std_logic;
signal heap_bh30_w81_11 :  std_logic;
signal heap_bh30_w80_10 :  std_logic;
signal heap_bh30_w79_11 :  std_logic;
signal heap_bh30_w78_11 :  std_logic;
signal heap_bh30_w77_10 :  std_logic;
signal heap_bh30_w76_11 :  std_logic;
signal heap_bh30_w75_11 :  std_logic;
signal heap_bh30_w74_10 :  std_logic;
signal heap_bh30_w73_11 :  std_logic;
signal heap_bh30_w72_11 :  std_logic;
signal heap_bh30_w71_10 :  std_logic;
signal heap_bh30_w70_10 :  std_logic;
signal heap_bh30_w69_10 :  std_logic;
signal heap_bh30_w68_9 :  std_logic;
signal heap_bh30_w67_10 :  std_logic;
signal heap_bh30_w66_9 :  std_logic;
signal heap_bh30_w65_8 :  std_logic;
signal heap_bh30_w64_9 :  std_logic;
signal heap_bh30_w63_8 :  std_logic;
signal heap_bh30_w62_7 :  std_logic;
signal heap_bh30_w61_8 :  std_logic;
signal heap_bh30_w60_8 :  std_logic;
signal heap_bh30_w59_7 :  std_logic;
signal heap_bh30_w58_8 :  std_logic;
signal heap_bh30_w57_8 :  std_logic;
signal heap_bh30_w56_7 :  std_logic;
signal heap_bh30_w55_8 :  std_logic;
signal heap_bh30_w54_8 :  std_logic;
signal heap_bh30_w53_7 :  std_logic;
signal heap_bh30_w52_8 :  std_logic;
signal heap_bh30_w51_8 :  std_logic;
signal heap_bh30_w50_7 :  std_logic;
signal heap_bh30_w49_7 :  std_logic;
signal heap_bh30_w48_7 :  std_logic;
signal heap_bh30_w47_6 :  std_logic;
signal DSP_bh30_ch18_0 :  std_logic_vector(40 downto 0);
signal heap_bh30_w63_9 :  std_logic;
signal heap_bh30_w62_8 :  std_logic;
signal heap_bh30_w61_9 :  std_logic;
signal heap_bh30_w60_9 :  std_logic;
signal heap_bh30_w59_8 :  std_logic;
signal heap_bh30_w58_9 :  std_logic;
signal heap_bh30_w57_9 :  std_logic;
signal heap_bh30_w56_8 :  std_logic;
signal heap_bh30_w55_9 :  std_logic;
signal heap_bh30_w54_9 :  std_logic;
signal heap_bh30_w53_8 :  std_logic;
signal heap_bh30_w52_9 :  std_logic;
signal heap_bh30_w51_9 :  std_logic;
signal heap_bh30_w50_8 :  std_logic;
signal heap_bh30_w49_8 :  std_logic;
signal heap_bh30_w48_8 :  std_logic;
signal heap_bh30_w47_7 :  std_logic;
signal heap_bh30_w46_7 :  std_logic;
signal heap_bh30_w45_7 :  std_logic;
signal heap_bh30_w44_6 :  std_logic;
signal heap_bh30_w43_7 :  std_logic;
signal heap_bh30_w42_7 :  std_logic;
signal heap_bh30_w41_6 :  std_logic;
signal heap_bh30_w40_7 :  std_logic;
signal heap_bh30_w39_6 :  std_logic;
signal heap_bh30_w38_5 :  std_logic;
signal heap_bh30_w37_6 :  std_logic;
signal heap_bh30_w36_6 :  std_logic;
signal heap_bh30_w35_5 :  std_logic;
signal heap_bh30_w34_6 :  std_logic;
signal heap_bh30_w33_6 :  std_logic;
signal heap_bh30_w32_4 :  std_logic;
signal heap_bh30_w31_5 :  std_logic;
signal heap_bh30_w30_5 :  std_logic;
signal heap_bh30_w29_4 :  std_logic;
signal heap_bh30_w28_5 :  std_logic;
signal heap_bh30_w27_5 :  std_logic;
signal heap_bh30_w26_4 :  std_logic;
signal heap_bh30_w25_5 :  std_logic;
signal heap_bh30_w24_5 :  std_logic;
signal heap_bh30_w23_4 :  std_logic;
signal DSP_bh30_ch19_0 :  std_logic_vector(40 downto 0);
signal heap_bh30_w39_7 :  std_logic;
signal heap_bh30_w38_6 :  std_logic;
signal heap_bh30_w37_7 :  std_logic;
signal heap_bh30_w36_7 :  std_logic;
signal heap_bh30_w35_6 :  std_logic;
signal heap_bh30_w34_7 :  std_logic;
signal heap_bh30_w33_7 :  std_logic;
signal heap_bh30_w32_5 :  std_logic;
signal heap_bh30_w31_6 :  std_logic;
signal heap_bh30_w30_6 :  std_logic;
signal heap_bh30_w29_5 :  std_logic;
signal heap_bh30_w28_6 :  std_logic;
signal heap_bh30_w27_6 :  std_logic;
signal heap_bh30_w26_5 :  std_logic;
signal heap_bh30_w25_6 :  std_logic;
signal heap_bh30_w24_6 :  std_logic;
signal heap_bh30_w23_5 :  std_logic;
signal heap_bh30_w22_5 :  std_logic;
signal heap_bh30_w21_5 :  std_logic;
signal heap_bh30_w20_4 :  std_logic;
signal heap_bh30_w19_5 :  std_logic;
signal heap_bh30_w18_5 :  std_logic;
signal heap_bh30_w17_4 :  std_logic;
signal heap_bh30_w16_5 :  std_logic;
signal heap_bh30_w15_4 :  std_logic;
signal heap_bh30_w14_3 :  std_logic;
signal heap_bh30_w13_4 :  std_logic;
signal heap_bh30_w12_4 :  std_logic;
signal heap_bh30_w11_3 :  std_logic;
signal heap_bh30_w10_4 :  std_logic;
signal heap_bh30_w9_4 :  std_logic;
signal heap_bh30_w8_3 :  std_logic;
signal heap_bh30_w7_4 :  std_logic;
signal heap_bh30_w6_4 :  std_logic;
signal heap_bh30_w5_3 :  std_logic;
signal heap_bh30_w4_3 :  std_logic;
signal heap_bh30_w3_3 :  std_logic;
signal heap_bh30_w2_2 :  std_logic;
signal heap_bh30_w1_1 :  std_logic;
signal heap_bh30_w0_1 :  std_logic;
signal CompressorIn_bh30_0_0 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_0_1 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_0_0 :  std_logic_vector(2 downto 0);
signal heap_bh30_w6_5 :  std_logic;
signal heap_bh30_w7_5 :  std_logic;
signal heap_bh30_w8_4 :  std_logic;
signal CompressorIn_bh30_1_2 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_1_3 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_1_1 :  std_logic_vector(2 downto 0);
signal heap_bh30_w9_5 :  std_logic;
signal heap_bh30_w10_5 :  std_logic;
signal heap_bh30_w11_4 :  std_logic;
signal CompressorIn_bh30_2_4 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_2_5 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_2_2 :  std_logic_vector(2 downto 0);
signal heap_bh30_w12_5 :  std_logic;
signal heap_bh30_w13_5 :  std_logic;
signal heap_bh30_w14_4 :  std_logic;
signal CompressorIn_bh30_3_6 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_3_7 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_3_3 :  std_logic_vector(2 downto 0);
signal heap_bh30_w15_5 :  std_logic;
signal heap_bh30_w16_6 :  std_logic;
signal heap_bh30_w17_5 :  std_logic;
signal CompressorIn_bh30_4_8 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_4_9 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_4_4 :  std_logic_vector(2 downto 0);
signal heap_bh30_w18_6 :  std_logic;
signal heap_bh30_w19_6 :  std_logic;
signal heap_bh30_w20_5 :  std_logic;
signal CompressorIn_bh30_5_10 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_5_11 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_5_5 :  std_logic_vector(2 downto 0);
signal heap_bh30_w21_6 :  std_logic;
signal heap_bh30_w22_6 :  std_logic;
signal heap_bh30_w23_6 :  std_logic;
signal CompressorIn_bh30_6_12 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_6_13 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_6_6 :  std_logic_vector(2 downto 0);
signal heap_bh30_w24_7 :  std_logic;
signal heap_bh30_w25_7 :  std_logic;
signal heap_bh30_w26_6 :  std_logic;
signal CompressorIn_bh30_7_14 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_7_15 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_7_7 :  std_logic_vector(2 downto 0);
signal heap_bh30_w27_7 :  std_logic;
signal heap_bh30_w28_7 :  std_logic;
signal heap_bh30_w29_6 :  std_logic;
signal CompressorIn_bh30_8_16 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_8_17 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_8_8 :  std_logic_vector(2 downto 0);
signal heap_bh30_w30_7 :  std_logic;
signal heap_bh30_w31_7 :  std_logic;
signal heap_bh30_w32_6 :  std_logic;
signal CompressorIn_bh30_9_18 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_9_19 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_9_9 :  std_logic_vector(2 downto 0);
signal heap_bh30_w33_8 :  std_logic;
signal heap_bh30_w34_8 :  std_logic;
signal heap_bh30_w35_7 :  std_logic;
signal CompressorIn_bh30_10_20 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_10_21 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_10_10 :  std_logic_vector(2 downto 0);
signal heap_bh30_w36_8 :  std_logic;
signal heap_bh30_w37_8 :  std_logic;
signal heap_bh30_w38_7 :  std_logic;
signal CompressorIn_bh30_11_22 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_11_23 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_11_11 :  std_logic_vector(2 downto 0);
signal heap_bh30_w39_8 :  std_logic;
signal heap_bh30_w40_8 :  std_logic;
signal heap_bh30_w41_7 :  std_logic;
signal CompressorIn_bh30_12_24 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_12_25 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_12_12 :  std_logic_vector(2 downto 0);
signal heap_bh30_w42_8 :  std_logic;
signal heap_bh30_w43_8 :  std_logic;
signal heap_bh30_w44_7 :  std_logic;
signal CompressorIn_bh30_13_26 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_13_27 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_13_13 :  std_logic_vector(2 downto 0);
signal heap_bh30_w45_8 :  std_logic;
signal heap_bh30_w46_8 :  std_logic;
signal heap_bh30_w47_8 :  std_logic;
signal CompressorIn_bh30_14_28 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_14_29 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_14_14 :  std_logic_vector(2 downto 0);
signal heap_bh30_w48_9 :  std_logic;
signal heap_bh30_w49_9 :  std_logic;
signal heap_bh30_w50_9 :  std_logic;
signal CompressorIn_bh30_15_30 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_15_31 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_15_15 :  std_logic_vector(2 downto 0);
signal heap_bh30_w51_10 :  std_logic;
signal heap_bh30_w52_10 :  std_logic;
signal heap_bh30_w53_9 :  std_logic;
signal CompressorIn_bh30_16_32 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_16_33 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_16_16 :  std_logic_vector(2 downto 0);
signal heap_bh30_w54_10 :  std_logic;
signal heap_bh30_w55_10 :  std_logic;
signal heap_bh30_w56_9 :  std_logic;
signal CompressorIn_bh30_17_34 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_17_35 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_17_17 :  std_logic_vector(2 downto 0);
signal heap_bh30_w57_10 :  std_logic;
signal heap_bh30_w58_10 :  std_logic;
signal heap_bh30_w59_9 :  std_logic;
signal CompressorIn_bh30_18_36 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_18_37 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_18_18 :  std_logic_vector(2 downto 0);
signal heap_bh30_w60_10 :  std_logic;
signal heap_bh30_w61_10 :  std_logic;
signal heap_bh30_w62_9 :  std_logic;
signal CompressorIn_bh30_19_38 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_19_39 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_19_19 :  std_logic_vector(2 downto 0);
signal heap_bh30_w63_10 :  std_logic;
signal heap_bh30_w64_10 :  std_logic;
signal heap_bh30_w65_9 :  std_logic;
signal CompressorIn_bh30_20_40 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_20_41 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_20_20 :  std_logic_vector(2 downto 0);
signal heap_bh30_w66_10 :  std_logic;
signal heap_bh30_w67_11 :  std_logic;
signal heap_bh30_w68_10 :  std_logic;
signal CompressorIn_bh30_21_42 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_21_43 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_21_21 :  std_logic_vector(2 downto 0);
signal heap_bh30_w69_11 :  std_logic;
signal heap_bh30_w70_11 :  std_logic;
signal heap_bh30_w71_11 :  std_logic;
signal CompressorIn_bh30_22_44 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_22_45 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_22_22 :  std_logic_vector(2 downto 0);
signal heap_bh30_w72_12 :  std_logic;
signal heap_bh30_w73_12 :  std_logic;
signal heap_bh30_w74_11 :  std_logic;
signal CompressorIn_bh30_23_46 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_23_47 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_23_23 :  std_logic_vector(2 downto 0);
signal heap_bh30_w75_12 :  std_logic;
signal heap_bh30_w76_12 :  std_logic;
signal heap_bh30_w77_11 :  std_logic;
signal CompressorIn_bh30_24_48 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_24_49 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_24_24 :  std_logic_vector(2 downto 0);
signal heap_bh30_w78_12 :  std_logic;
signal heap_bh30_w79_12 :  std_logic;
signal heap_bh30_w80_11 :  std_logic;
signal CompressorIn_bh30_25_50 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_25_51 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_25_25 :  std_logic_vector(2 downto 0);
signal heap_bh30_w81_12 :  std_logic;
signal heap_bh30_w82_12 :  std_logic;
signal heap_bh30_w83_11 :  std_logic;
signal CompressorIn_bh30_26_52 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_26_53 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_26_26 :  std_logic_vector(2 downto 0);
signal heap_bh30_w84_12 :  std_logic;
signal heap_bh30_w85_12 :  std_logic;
signal heap_bh30_w86_11 :  std_logic;
signal CompressorIn_bh30_27_54 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_27_55 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_27_27 :  std_logic_vector(2 downto 0);
signal heap_bh30_w87_12 :  std_logic;
signal heap_bh30_w88_12 :  std_logic;
signal heap_bh30_w89_11 :  std_logic;
signal CompressorIn_bh30_28_56 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_28_57 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_28_28 :  std_logic_vector(2 downto 0);
signal heap_bh30_w3_4 :  std_logic;
signal heap_bh30_w4_4 :  std_logic;
signal heap_bh30_w5_4 :  std_logic;
signal CompressorIn_bh30_29_58 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_29_59 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_29_29 :  std_logic_vector(2 downto 0);
signal heap_bh30_w7_6 :  std_logic;
signal heap_bh30_w8_5 :  std_logic;
signal heap_bh30_w9_6 :  std_logic;
signal CompressorIn_bh30_30_60 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_30_61 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_30_30 :  std_logic_vector(2 downto 0);
signal heap_bh30_w10_6 :  std_logic;
signal heap_bh30_w11_5 :  std_logic;
signal heap_bh30_w12_6 :  std_logic;
signal CompressorIn_bh30_31_62 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_31_63 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_31_31 :  std_logic_vector(2 downto 0);
signal heap_bh30_w13_6 :  std_logic;
signal heap_bh30_w14_5 :  std_logic;
signal heap_bh30_w15_6 :  std_logic;
signal CompressorIn_bh30_32_64 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_32_65 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_32_32 :  std_logic_vector(2 downto 0);
signal heap_bh30_w16_7 :  std_logic;
signal heap_bh30_w17_6 :  std_logic;
signal heap_bh30_w18_7 :  std_logic;
signal CompressorIn_bh30_33_66 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_33_67 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_33_33 :  std_logic_vector(2 downto 0);
signal heap_bh30_w19_7 :  std_logic;
signal heap_bh30_w20_6 :  std_logic;
signal heap_bh30_w21_7 :  std_logic;
signal CompressorIn_bh30_34_68 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_34_69 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_34_34 :  std_logic_vector(2 downto 0);
signal heap_bh30_w22_7 :  std_logic;
signal heap_bh30_w23_7 :  std_logic;
signal heap_bh30_w24_8 :  std_logic;
signal CompressorIn_bh30_35_70 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_35_71 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_35_35 :  std_logic_vector(2 downto 0);
signal heap_bh30_w25_8 :  std_logic;
signal heap_bh30_w26_7 :  std_logic;
signal heap_bh30_w27_8 :  std_logic;
signal CompressorIn_bh30_36_72 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_36_73 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_36_36 :  std_logic_vector(2 downto 0);
signal heap_bh30_w28_8 :  std_logic;
signal heap_bh30_w29_7 :  std_logic;
signal heap_bh30_w30_8 :  std_logic;
signal CompressorIn_bh30_37_74 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_37_75 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_37_37 :  std_logic_vector(2 downto 0);
signal heap_bh30_w31_8 :  std_logic;
signal heap_bh30_w32_7 :  std_logic;
signal heap_bh30_w33_9 :  std_logic;
signal CompressorIn_bh30_38_76 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_38_77 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_38_38 :  std_logic_vector(2 downto 0);
signal heap_bh30_w34_9 :  std_logic;
signal heap_bh30_w35_8 :  std_logic;
signal heap_bh30_w36_9 :  std_logic;
signal CompressorIn_bh30_39_78 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_39_79 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_39_39 :  std_logic_vector(2 downto 0);
signal heap_bh30_w37_9 :  std_logic;
signal heap_bh30_w38_8 :  std_logic;
signal heap_bh30_w39_9 :  std_logic;
signal CompressorIn_bh30_40_80 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_40_81 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_40_40 :  std_logic_vector(2 downto 0);
signal heap_bh30_w40_9 :  std_logic;
signal heap_bh30_w41_8 :  std_logic;
signal heap_bh30_w42_9 :  std_logic;
signal CompressorIn_bh30_41_82 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_41_83 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_41_41 :  std_logic_vector(2 downto 0);
signal heap_bh30_w43_9 :  std_logic;
signal heap_bh30_w44_8 :  std_logic;
signal heap_bh30_w45_9 :  std_logic;
signal CompressorIn_bh30_42_84 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_42_85 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_42_42 :  std_logic_vector(2 downto 0);
signal heap_bh30_w46_9 :  std_logic;
signal heap_bh30_w47_9 :  std_logic;
signal heap_bh30_w48_10 :  std_logic;
signal CompressorIn_bh30_43_86 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_43_87 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_43_43 :  std_logic_vector(2 downto 0);
signal heap_bh30_w49_10 :  std_logic;
signal heap_bh30_w50_10 :  std_logic;
signal heap_bh30_w51_11 :  std_logic;
signal CompressorIn_bh30_44_88 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_44_89 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_44_44 :  std_logic_vector(2 downto 0);
signal heap_bh30_w52_11 :  std_logic;
signal heap_bh30_w53_10 :  std_logic;
signal heap_bh30_w54_11 :  std_logic;
signal CompressorIn_bh30_45_90 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_45_91 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_45_45 :  std_logic_vector(2 downto 0);
signal heap_bh30_w55_11 :  std_logic;
signal heap_bh30_w56_10 :  std_logic;
signal heap_bh30_w57_11 :  std_logic;
signal CompressorIn_bh30_46_92 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_46_93 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_46_46 :  std_logic_vector(2 downto 0);
signal heap_bh30_w58_11 :  std_logic;
signal heap_bh30_w59_10 :  std_logic;
signal heap_bh30_w60_11 :  std_logic;
signal CompressorIn_bh30_47_94 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_47_95 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_47_47 :  std_logic_vector(2 downto 0);
signal heap_bh30_w61_11 :  std_logic;
signal heap_bh30_w62_10 :  std_logic;
signal heap_bh30_w63_11 :  std_logic;
signal CompressorIn_bh30_48_96 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_48_97 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_48_48 :  std_logic_vector(2 downto 0);
signal heap_bh30_w64_11 :  std_logic;
signal heap_bh30_w65_10 :  std_logic;
signal heap_bh30_w66_11 :  std_logic;
signal CompressorIn_bh30_49_98 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_49_99 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_49_49 :  std_logic_vector(2 downto 0);
signal heap_bh30_w67_12 :  std_logic;
signal heap_bh30_w68_11 :  std_logic;
signal heap_bh30_w69_12 :  std_logic;
signal CompressorIn_bh30_50_100 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_50_101 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_50_50 :  std_logic_vector(2 downto 0);
signal heap_bh30_w70_12 :  std_logic;
signal heap_bh30_w71_12 :  std_logic;
signal heap_bh30_w72_13 :  std_logic;
signal CompressorIn_bh30_51_102 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_51_103 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_51_51 :  std_logic_vector(2 downto 0);
signal heap_bh30_w73_13 :  std_logic;
signal heap_bh30_w74_12 :  std_logic;
signal heap_bh30_w75_13 :  std_logic;
signal CompressorIn_bh30_52_104 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_52_105 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_52_52 :  std_logic_vector(2 downto 0);
signal heap_bh30_w76_13 :  std_logic;
signal heap_bh30_w77_12 :  std_logic;
signal heap_bh30_w78_13 :  std_logic;
signal CompressorIn_bh30_53_106 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_53_107 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_53_53 :  std_logic_vector(2 downto 0);
signal heap_bh30_w79_13 :  std_logic;
signal heap_bh30_w80_12 :  std_logic;
signal heap_bh30_w81_13 :  std_logic;
signal CompressorIn_bh30_54_108 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_54_109 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_54_54 :  std_logic_vector(2 downto 0);
signal heap_bh30_w82_13 :  std_logic;
signal heap_bh30_w83_12 :  std_logic;
signal heap_bh30_w84_13 :  std_logic;
signal CompressorIn_bh30_55_110 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_55_111 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_55_55 :  std_logic_vector(2 downto 0);
signal heap_bh30_w85_13 :  std_logic;
signal heap_bh30_w86_12 :  std_logic;
signal heap_bh30_w87_13 :  std_logic;
signal CompressorIn_bh30_56_112 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_56_113 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_56_56 :  std_logic_vector(2 downto 0);
signal heap_bh30_w88_13 :  std_logic;
signal heap_bh30_w89_12 :  std_logic;
signal heap_bh30_w90_11 :  std_logic;
signal CompressorIn_bh30_57_114 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_57_115 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_57_57 :  std_logic_vector(2 downto 0);
signal heap_bh30_w90_12 :  std_logic;
signal heap_bh30_w91_11 :  std_logic;
signal heap_bh30_w92_9 :  std_logic;
signal CompressorIn_bh30_58_116 :  std_logic_vector(2 downto 0);
signal CompressorOut_bh30_58_58 :  std_logic_vector(1 downto 0);
signal heap_bh30_w5_5 :  std_logic;
signal heap_bh30_w6_6 :  std_logic;
signal CompressorIn_bh30_59_117 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_59_118 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_59_59 :  std_logic_vector(2 downto 0);
signal heap_bh30_w8_6 :  std_logic;
signal heap_bh30_w9_7 :  std_logic;
signal heap_bh30_w10_7 :  std_logic;
signal CompressorIn_bh30_60_119 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_60_120 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_60_60 :  std_logic_vector(2 downto 0);
signal heap_bh30_w11_6 :  std_logic;
signal heap_bh30_w12_7 :  std_logic;
signal heap_bh30_w13_7 :  std_logic;
signal CompressorIn_bh30_61_121 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_61_122 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_61_61 :  std_logic_vector(2 downto 0);
signal heap_bh30_w14_6 :  std_logic;
signal heap_bh30_w15_7 :  std_logic;
signal heap_bh30_w16_8 :  std_logic;
signal CompressorIn_bh30_62_123 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_62_124 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_62_62 :  std_logic_vector(2 downto 0);
signal heap_bh30_w17_7 :  std_logic;
signal heap_bh30_w18_8 :  std_logic;
signal heap_bh30_w19_8 :  std_logic;
signal CompressorIn_bh30_63_125 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_63_126 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_63_63 :  std_logic_vector(2 downto 0);
signal heap_bh30_w20_7 :  std_logic;
signal heap_bh30_w21_8 :  std_logic;
signal heap_bh30_w22_8 :  std_logic;
signal CompressorIn_bh30_64_127 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_64_128 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_64_64 :  std_logic_vector(2 downto 0);
signal heap_bh30_w23_8 :  std_logic;
signal heap_bh30_w24_9 :  std_logic;
signal heap_bh30_w25_9 :  std_logic;
signal CompressorIn_bh30_65_129 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_65_130 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_65_65 :  std_logic_vector(2 downto 0);
signal heap_bh30_w26_8 :  std_logic;
signal heap_bh30_w27_9 :  std_logic;
signal heap_bh30_w28_9 :  std_logic;
signal CompressorIn_bh30_66_131 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_66_132 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_66_66 :  std_logic_vector(2 downto 0);
signal heap_bh30_w29_8 :  std_logic;
signal heap_bh30_w30_9 :  std_logic;
signal heap_bh30_w31_9 :  std_logic;
signal CompressorIn_bh30_67_133 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_67_134 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_67_67 :  std_logic_vector(2 downto 0);
signal heap_bh30_w32_8 :  std_logic;
signal heap_bh30_w33_10 :  std_logic;
signal heap_bh30_w34_10 :  std_logic;
signal CompressorIn_bh30_68_135 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_68_136 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_68_68 :  std_logic_vector(2 downto 0);
signal heap_bh30_w35_9 :  std_logic;
signal heap_bh30_w36_10 :  std_logic;
signal heap_bh30_w37_10 :  std_logic;
signal CompressorIn_bh30_69_137 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_69_138 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_69_69 :  std_logic_vector(2 downto 0);
signal heap_bh30_w38_9 :  std_logic;
signal heap_bh30_w39_10 :  std_logic;
signal heap_bh30_w40_10 :  std_logic;
signal CompressorIn_bh30_70_139 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_70_140 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_70_70 :  std_logic_vector(2 downto 0);
signal heap_bh30_w41_9 :  std_logic;
signal heap_bh30_w42_10 :  std_logic;
signal heap_bh30_w43_10 :  std_logic;
signal CompressorIn_bh30_71_141 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_71_142 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_71_71 :  std_logic_vector(2 downto 0);
signal heap_bh30_w44_9 :  std_logic;
signal heap_bh30_w45_10 :  std_logic;
signal heap_bh30_w46_10 :  std_logic;
signal CompressorIn_bh30_72_143 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_72_144 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_72_72 :  std_logic_vector(2 downto 0);
signal heap_bh30_w47_10 :  std_logic;
signal heap_bh30_w48_11 :  std_logic;
signal heap_bh30_w49_11 :  std_logic;
signal CompressorIn_bh30_73_145 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_73_146 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_73_73 :  std_logic_vector(2 downto 0);
signal heap_bh30_w50_11 :  std_logic;
signal heap_bh30_w51_12 :  std_logic;
signal heap_bh30_w52_12 :  std_logic;
signal CompressorIn_bh30_74_147 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_74_148 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_74_74 :  std_logic_vector(2 downto 0);
signal heap_bh30_w53_11 :  std_logic;
signal heap_bh30_w54_12 :  std_logic;
signal heap_bh30_w55_12 :  std_logic;
signal CompressorIn_bh30_75_149 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_75_150 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_75_75 :  std_logic_vector(2 downto 0);
signal heap_bh30_w56_11 :  std_logic;
signal heap_bh30_w57_12 :  std_logic;
signal heap_bh30_w58_12 :  std_logic;
signal CompressorIn_bh30_76_151 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_76_152 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_76_76 :  std_logic_vector(2 downto 0);
signal heap_bh30_w59_11 :  std_logic;
signal heap_bh30_w60_12 :  std_logic;
signal heap_bh30_w61_12 :  std_logic;
signal CompressorIn_bh30_77_153 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_77_154 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_77_77 :  std_logic_vector(2 downto 0);
signal heap_bh30_w62_11 :  std_logic;
signal heap_bh30_w63_12 :  std_logic;
signal heap_bh30_w64_12 :  std_logic;
signal CompressorIn_bh30_78_155 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_78_156 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_78_78 :  std_logic_vector(2 downto 0);
signal heap_bh30_w65_11 :  std_logic;
signal heap_bh30_w66_12 :  std_logic;
signal heap_bh30_w67_13 :  std_logic;
signal CompressorIn_bh30_79_157 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_79_158 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_79_79 :  std_logic_vector(2 downto 0);
signal heap_bh30_w68_12 :  std_logic;
signal heap_bh30_w69_13 :  std_logic;
signal heap_bh30_w70_13 :  std_logic;
signal CompressorIn_bh30_80_159 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_80_160 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_80_80 :  std_logic_vector(2 downto 0);
signal heap_bh30_w71_13 :  std_logic;
signal heap_bh30_w72_14 :  std_logic;
signal heap_bh30_w73_14 :  std_logic;
signal CompressorIn_bh30_81_161 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_81_162 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_81_81 :  std_logic_vector(2 downto 0);
signal heap_bh30_w74_13 :  std_logic;
signal heap_bh30_w75_14 :  std_logic;
signal heap_bh30_w76_14 :  std_logic;
signal CompressorIn_bh30_82_163 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_82_164 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_82_82 :  std_logic_vector(2 downto 0);
signal heap_bh30_w77_13 :  std_logic;
signal heap_bh30_w78_14 :  std_logic;
signal heap_bh30_w79_14 :  std_logic;
signal CompressorIn_bh30_83_165 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_83_166 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_83_83 :  std_logic_vector(2 downto 0);
signal heap_bh30_w80_13 :  std_logic;
signal heap_bh30_w81_14 :  std_logic;
signal heap_bh30_w82_14 :  std_logic;
signal CompressorIn_bh30_84_167 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_84_168 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_84_84 :  std_logic_vector(2 downto 0);
signal heap_bh30_w83_13 :  std_logic;
signal heap_bh30_w84_14 :  std_logic;
signal heap_bh30_w85_14 :  std_logic;
signal CompressorIn_bh30_85_169 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_85_170 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_85_85 :  std_logic_vector(2 downto 0);
signal heap_bh30_w86_13 :  std_logic;
signal heap_bh30_w87_14 :  std_logic;
signal heap_bh30_w88_14 :  std_logic;
signal CompressorIn_bh30_86_171 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_86_172 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_86_86 :  std_logic_vector(2 downto 0);
signal heap_bh30_w89_13 :  std_logic;
signal heap_bh30_w90_13 :  std_logic;
signal heap_bh30_w91_12 :  std_logic;
signal CompressorIn_bh30_87_173 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_87_174 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_87_87 :  std_logic_vector(2 downto 0);
signal heap_bh30_w91_13 :  std_logic;
signal heap_bh30_w92_10 :  std_logic;
signal heap_bh30_w93_9 :  std_logic;
signal CompressorIn_bh30_88_175 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_88_176 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_88_88 :  std_logic_vector(2 downto 0);
signal heap_bh30_w10_8 :  std_logic;
signal heap_bh30_w11_7 :  std_logic;
signal heap_bh30_w12_8 :  std_logic;
signal CompressorIn_bh30_89_177 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_89_178 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_89_89 :  std_logic_vector(2 downto 0);
signal heap_bh30_w13_8 :  std_logic;
signal heap_bh30_w14_7 :  std_logic;
signal heap_bh30_w15_8 :  std_logic;
signal CompressorIn_bh30_90_179 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_90_180 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_90_90 :  std_logic_vector(2 downto 0);
signal heap_bh30_w16_9 :  std_logic;
signal heap_bh30_w17_8 :  std_logic;
signal heap_bh30_w18_9 :  std_logic;
signal CompressorIn_bh30_91_181 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_91_182 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_91_91 :  std_logic_vector(2 downto 0);
signal heap_bh30_w19_9 :  std_logic;
signal heap_bh30_w20_8 :  std_logic;
signal heap_bh30_w21_9 :  std_logic;
signal CompressorIn_bh30_92_183 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_92_184 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_92_92 :  std_logic_vector(2 downto 0);
signal heap_bh30_w22_9 :  std_logic;
signal heap_bh30_w23_9 :  std_logic;
signal heap_bh30_w24_10 :  std_logic;
signal CompressorIn_bh30_93_185 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_93_186 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_93_93 :  std_logic_vector(2 downto 0);
signal heap_bh30_w25_10 :  std_logic;
signal heap_bh30_w26_9 :  std_logic;
signal heap_bh30_w27_10 :  std_logic;
signal CompressorIn_bh30_94_187 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_94_188 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_94_94 :  std_logic_vector(2 downto 0);
signal heap_bh30_w28_10 :  std_logic;
signal heap_bh30_w29_9 :  std_logic;
signal heap_bh30_w30_10 :  std_logic;
signal CompressorIn_bh30_95_189 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_95_190 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_95_95 :  std_logic_vector(2 downto 0);
signal heap_bh30_w31_10 :  std_logic;
signal heap_bh30_w32_9 :  std_logic;
signal heap_bh30_w33_11 :  std_logic;
signal CompressorIn_bh30_96_191 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_96_192 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_96_96 :  std_logic_vector(2 downto 0);
signal heap_bh30_w34_11 :  std_logic;
signal heap_bh30_w35_10 :  std_logic;
signal heap_bh30_w36_11 :  std_logic;
signal CompressorIn_bh30_97_193 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_97_194 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_97_97 :  std_logic_vector(2 downto 0);
signal heap_bh30_w37_11 :  std_logic;
signal heap_bh30_w38_10 :  std_logic;
signal heap_bh30_w39_11 :  std_logic;
signal CompressorIn_bh30_98_195 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_98_196 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_98_98 :  std_logic_vector(2 downto 0);
signal heap_bh30_w40_11 :  std_logic;
signal heap_bh30_w41_10 :  std_logic;
signal heap_bh30_w42_11 :  std_logic;
signal CompressorIn_bh30_99_197 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_99_198 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_99_99 :  std_logic_vector(2 downto 0);
signal heap_bh30_w43_11 :  std_logic;
signal heap_bh30_w44_10 :  std_logic;
signal heap_bh30_w45_11 :  std_logic;
signal CompressorIn_bh30_100_199 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_100_200 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_100_100 :  std_logic_vector(2 downto 0);
signal heap_bh30_w46_11 :  std_logic;
signal heap_bh30_w47_11 :  std_logic;
signal heap_bh30_w48_12 :  std_logic;
signal CompressorIn_bh30_101_201 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_101_202 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_101_101 :  std_logic_vector(2 downto 0);
signal heap_bh30_w49_12 :  std_logic;
signal heap_bh30_w50_12 :  std_logic;
signal heap_bh30_w51_13 :  std_logic;
signal CompressorIn_bh30_102_203 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_102_204 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_102_102 :  std_logic_vector(2 downto 0);
signal heap_bh30_w52_13 :  std_logic;
signal heap_bh30_w53_12 :  std_logic;
signal heap_bh30_w54_13 :  std_logic;
signal CompressorIn_bh30_103_205 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_103_206 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_103_103 :  std_logic_vector(2 downto 0);
signal heap_bh30_w55_13 :  std_logic;
signal heap_bh30_w56_12 :  std_logic;
signal heap_bh30_w57_13 :  std_logic;
signal CompressorIn_bh30_104_207 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_104_208 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_104_104 :  std_logic_vector(2 downto 0);
signal heap_bh30_w58_13 :  std_logic;
signal heap_bh30_w59_12 :  std_logic;
signal heap_bh30_w60_13 :  std_logic;
signal CompressorIn_bh30_105_209 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_105_210 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_105_105 :  std_logic_vector(2 downto 0);
signal heap_bh30_w61_13 :  std_logic;
signal heap_bh30_w62_12 :  std_logic;
signal heap_bh30_w63_13 :  std_logic;
signal CompressorIn_bh30_106_211 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_106_212 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_106_106 :  std_logic_vector(2 downto 0);
signal heap_bh30_w64_13 :  std_logic;
signal heap_bh30_w65_12 :  std_logic;
signal heap_bh30_w66_13 :  std_logic;
signal CompressorIn_bh30_107_213 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_107_214 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_107_107 :  std_logic_vector(2 downto 0);
signal heap_bh30_w67_14 :  std_logic;
signal heap_bh30_w68_13 :  std_logic;
signal heap_bh30_w69_14 :  std_logic;
signal CompressorIn_bh30_108_215 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_108_216 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_108_108 :  std_logic_vector(2 downto 0);
signal heap_bh30_w70_14 :  std_logic;
signal heap_bh30_w71_14 :  std_logic;
signal heap_bh30_w72_15 :  std_logic;
signal CompressorIn_bh30_109_217 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_109_218 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_109_109 :  std_logic_vector(2 downto 0);
signal heap_bh30_w73_15 :  std_logic;
signal heap_bh30_w74_14 :  std_logic;
signal heap_bh30_w75_15 :  std_logic;
signal CompressorIn_bh30_110_219 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_110_220 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_110_110 :  std_logic_vector(2 downto 0);
signal heap_bh30_w76_15 :  std_logic;
signal heap_bh30_w77_14 :  std_logic;
signal heap_bh30_w78_15 :  std_logic;
signal CompressorIn_bh30_111_221 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_111_222 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_111_111 :  std_logic_vector(2 downto 0);
signal heap_bh30_w79_15 :  std_logic;
signal heap_bh30_w80_14 :  std_logic;
signal heap_bh30_w81_15 :  std_logic;
signal CompressorIn_bh30_112_223 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_112_224 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_112_112 :  std_logic_vector(2 downto 0);
signal heap_bh30_w82_15 :  std_logic;
signal heap_bh30_w83_14 :  std_logic;
signal heap_bh30_w84_15 :  std_logic;
signal CompressorIn_bh30_113_225 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_113_226 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_113_113 :  std_logic_vector(2 downto 0);
signal heap_bh30_w85_15 :  std_logic;
signal heap_bh30_w86_14 :  std_logic;
signal heap_bh30_w87_15 :  std_logic;
signal CompressorIn_bh30_114_227 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_114_228 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_114_114 :  std_logic_vector(2 downto 0);
signal heap_bh30_w88_15 :  std_logic;
signal heap_bh30_w89_14 :  std_logic;
signal heap_bh30_w90_14 :  std_logic;
signal CompressorIn_bh30_115_229 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_115_115 :  std_logic_vector(2 downto 0);
signal heap_bh30_w33_12 :  std_logic;
signal heap_bh30_w34_12 :  std_logic;
signal heap_bh30_w35_11 :  std_logic;
signal CompressorIn_bh30_116_230 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_116_116 :  std_logic_vector(2 downto 0);
signal heap_bh30_w36_12 :  std_logic;
signal heap_bh30_w37_12 :  std_logic;
signal heap_bh30_w38_11 :  std_logic;
signal CompressorIn_bh30_117_231 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_117_117 :  std_logic_vector(2 downto 0);
signal heap_bh30_w39_12 :  std_logic;
signal heap_bh30_w40_12 :  std_logic;
signal heap_bh30_w41_11 :  std_logic;
signal CompressorIn_bh30_118_232 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_118_118 :  std_logic_vector(2 downto 0);
signal heap_bh30_w42_12 :  std_logic;
signal heap_bh30_w43_12 :  std_logic;
signal heap_bh30_w44_11 :  std_logic;
signal CompressorIn_bh30_119_233 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_119_119 :  std_logic_vector(2 downto 0);
signal heap_bh30_w45_12 :  std_logic;
signal heap_bh30_w46_12 :  std_logic;
signal heap_bh30_w47_12 :  std_logic;
signal CompressorIn_bh30_120_234 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_120_120 :  std_logic_vector(2 downto 0);
signal heap_bh30_w47_13 :  std_logic;
signal heap_bh30_w48_13 :  std_logic;
signal heap_bh30_w49_13 :  std_logic;
signal CompressorIn_bh30_121_235 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_121_121 :  std_logic_vector(2 downto 0);
signal heap_bh30_w48_14 :  std_logic;
signal heap_bh30_w49_14 :  std_logic;
signal heap_bh30_w50_13 :  std_logic;
signal CompressorIn_bh30_122_236 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_122_122 :  std_logic_vector(2 downto 0);
signal heap_bh30_w49_15 :  std_logic;
signal heap_bh30_w50_14 :  std_logic;
signal heap_bh30_w51_14 :  std_logic;
signal CompressorIn_bh30_123_237 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_123_123 :  std_logic_vector(2 downto 0);
signal heap_bh30_w50_15 :  std_logic;
signal heap_bh30_w51_15 :  std_logic;
signal heap_bh30_w52_14 :  std_logic;
signal CompressorIn_bh30_124_238 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_124_124 :  std_logic_vector(2 downto 0);
signal heap_bh30_w51_16 :  std_logic;
signal heap_bh30_w52_15 :  std_logic;
signal heap_bh30_w53_13 :  std_logic;
signal CompressorIn_bh30_125_239 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_125_125 :  std_logic_vector(2 downto 0);
signal heap_bh30_w52_16 :  std_logic;
signal heap_bh30_w53_14 :  std_logic;
signal heap_bh30_w54_14 :  std_logic;
signal CompressorIn_bh30_126_240 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_126_126 :  std_logic_vector(2 downto 0);
signal heap_bh30_w53_15 :  std_logic;
signal heap_bh30_w54_15 :  std_logic;
signal heap_bh30_w55_14 :  std_logic;
signal CompressorIn_bh30_127_241 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_127_127 :  std_logic_vector(2 downto 0);
signal heap_bh30_w54_16 :  std_logic;
signal heap_bh30_w55_15 :  std_logic;
signal heap_bh30_w56_13 :  std_logic;
signal CompressorIn_bh30_128_242 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_128_128 :  std_logic_vector(2 downto 0);
signal heap_bh30_w55_16 :  std_logic;
signal heap_bh30_w56_14 :  std_logic;
signal heap_bh30_w57_14 :  std_logic;
signal CompressorIn_bh30_129_243 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_129_129 :  std_logic_vector(2 downto 0);
signal heap_bh30_w56_15 :  std_logic;
signal heap_bh30_w57_15 :  std_logic;
signal heap_bh30_w58_14 :  std_logic;
signal CompressorIn_bh30_130_244 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_130_130 :  std_logic_vector(2 downto 0);
signal heap_bh30_w57_16 :  std_logic;
signal heap_bh30_w58_15 :  std_logic;
signal heap_bh30_w59_13 :  std_logic;
signal CompressorIn_bh30_131_245 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_131_131 :  std_logic_vector(2 downto 0);
signal heap_bh30_w58_16 :  std_logic;
signal heap_bh30_w59_14 :  std_logic;
signal heap_bh30_w60_14 :  std_logic;
signal CompressorIn_bh30_132_246 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_132_132 :  std_logic_vector(2 downto 0);
signal heap_bh30_w59_15 :  std_logic;
signal heap_bh30_w60_15 :  std_logic;
signal heap_bh30_w61_14 :  std_logic;
signal CompressorIn_bh30_133_247 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_133_133 :  std_logic_vector(2 downto 0);
signal heap_bh30_w60_16 :  std_logic;
signal heap_bh30_w61_15 :  std_logic;
signal heap_bh30_w62_13 :  std_logic;
signal CompressorIn_bh30_134_248 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_134_134 :  std_logic_vector(2 downto 0);
signal heap_bh30_w61_16 :  std_logic;
signal heap_bh30_w62_14 :  std_logic;
signal heap_bh30_w63_14 :  std_logic;
signal CompressorIn_bh30_135_249 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_135_135 :  std_logic_vector(2 downto 0);
signal heap_bh30_w62_15 :  std_logic;
signal heap_bh30_w63_15 :  std_logic;
signal heap_bh30_w64_14 :  std_logic;
signal CompressorIn_bh30_136_250 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_136_136 :  std_logic_vector(2 downto 0);
signal heap_bh30_w63_16 :  std_logic;
signal heap_bh30_w64_15 :  std_logic;
signal heap_bh30_w65_13 :  std_logic;
signal CompressorIn_bh30_137_251 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_137_137 :  std_logic_vector(2 downto 0);
signal heap_bh30_w64_16 :  std_logic;
signal heap_bh30_w65_14 :  std_logic;
signal heap_bh30_w66_14 :  std_logic;
signal CompressorIn_bh30_138_252 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_138_138 :  std_logic_vector(2 downto 0);
signal heap_bh30_w65_15 :  std_logic;
signal heap_bh30_w66_15 :  std_logic;
signal heap_bh30_w67_15 :  std_logic;
signal CompressorIn_bh30_139_253 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_139_139 :  std_logic_vector(2 downto 0);
signal heap_bh30_w66_16 :  std_logic;
signal heap_bh30_w67_16 :  std_logic;
signal heap_bh30_w68_14 :  std_logic;
signal CompressorIn_bh30_140_254 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_140_140 :  std_logic_vector(2 downto 0);
signal heap_bh30_w67_17 :  std_logic;
signal heap_bh30_w68_15 :  std_logic;
signal heap_bh30_w69_15 :  std_logic;
signal CompressorIn_bh30_141_255 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_141_141 :  std_logic_vector(2 downto 0);
signal heap_bh30_w68_16 :  std_logic;
signal heap_bh30_w69_16 :  std_logic;
signal heap_bh30_w70_15 :  std_logic;
signal CompressorIn_bh30_142_256 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_142_142 :  std_logic_vector(2 downto 0);
signal heap_bh30_w69_17 :  std_logic;
signal heap_bh30_w70_16 :  std_logic;
signal heap_bh30_w71_15 :  std_logic;
signal CompressorIn_bh30_143_257 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_143_143 :  std_logic_vector(2 downto 0);
signal heap_bh30_w70_17 :  std_logic;
signal heap_bh30_w71_16 :  std_logic;
signal heap_bh30_w72_16 :  std_logic;
signal CompressorIn_bh30_144_258 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_144_144 :  std_logic_vector(2 downto 0);
signal heap_bh30_w71_17 :  std_logic;
signal heap_bh30_w72_17 :  std_logic;
signal heap_bh30_w73_16 :  std_logic;
signal CompressorIn_bh30_145_259 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_145_145 :  std_logic_vector(2 downto 0);
signal heap_bh30_w72_18 :  std_logic;
signal heap_bh30_w73_17 :  std_logic;
signal heap_bh30_w74_15 :  std_logic;
signal CompressorIn_bh30_146_260 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_146_146 :  std_logic_vector(2 downto 0);
signal heap_bh30_w73_18 :  std_logic;
signal heap_bh30_w74_16 :  std_logic;
signal heap_bh30_w75_16 :  std_logic;
signal CompressorIn_bh30_147_261 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_147_147 :  std_logic_vector(2 downto 0);
signal heap_bh30_w74_17 :  std_logic;
signal heap_bh30_w75_17 :  std_logic;
signal heap_bh30_w76_16 :  std_logic;
signal CompressorIn_bh30_148_262 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_148_148 :  std_logic_vector(2 downto 0);
signal heap_bh30_w75_18 :  std_logic;
signal heap_bh30_w76_17 :  std_logic;
signal heap_bh30_w77_15 :  std_logic;
signal CompressorIn_bh30_149_263 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_149_149 :  std_logic_vector(2 downto 0);
signal heap_bh30_w76_18 :  std_logic;
signal heap_bh30_w77_16 :  std_logic;
signal heap_bh30_w78_16 :  std_logic;
signal CompressorIn_bh30_150_264 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_150_150 :  std_logic_vector(2 downto 0);
signal heap_bh30_w77_17 :  std_logic;
signal heap_bh30_w78_17 :  std_logic;
signal heap_bh30_w79_16 :  std_logic;
signal CompressorIn_bh30_151_265 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_151_151 :  std_logic_vector(2 downto 0);
signal heap_bh30_w78_18 :  std_logic;
signal heap_bh30_w79_17 :  std_logic;
signal heap_bh30_w80_15 :  std_logic;
signal CompressorIn_bh30_152_266 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_152_152 :  std_logic_vector(2 downto 0);
signal heap_bh30_w79_18 :  std_logic;
signal heap_bh30_w80_16 :  std_logic;
signal heap_bh30_w81_16 :  std_logic;
signal CompressorIn_bh30_153_267 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_153_153 :  std_logic_vector(2 downto 0);
signal heap_bh30_w80_17 :  std_logic;
signal heap_bh30_w81_17 :  std_logic;
signal heap_bh30_w82_16 :  std_logic;
signal CompressorIn_bh30_154_268 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_154_154 :  std_logic_vector(2 downto 0);
signal heap_bh30_w81_18 :  std_logic;
signal heap_bh30_w82_17 :  std_logic;
signal heap_bh30_w83_15 :  std_logic;
signal CompressorIn_bh30_155_269 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_155_155 :  std_logic_vector(2 downto 0);
signal heap_bh30_w82_18 :  std_logic;
signal heap_bh30_w83_16 :  std_logic;
signal heap_bh30_w84_16 :  std_logic;
signal CompressorIn_bh30_156_270 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_156_156 :  std_logic_vector(2 downto 0);
signal heap_bh30_w83_17 :  std_logic;
signal heap_bh30_w84_17 :  std_logic;
signal heap_bh30_w85_16 :  std_logic;
signal CompressorIn_bh30_157_271 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_157_157 :  std_logic_vector(2 downto 0);
signal heap_bh30_w84_18 :  std_logic;
signal heap_bh30_w85_17 :  std_logic;
signal heap_bh30_w86_15 :  std_logic;
signal CompressorIn_bh30_158_272 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_158_158 :  std_logic_vector(2 downto 0);
signal heap_bh30_w85_18 :  std_logic;
signal heap_bh30_w86_16 :  std_logic;
signal heap_bh30_w87_16 :  std_logic;
signal CompressorIn_bh30_159_273 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_159_159 :  std_logic_vector(2 downto 0);
signal heap_bh30_w86_17 :  std_logic;
signal heap_bh30_w87_17 :  std_logic;
signal heap_bh30_w88_16 :  std_logic;
signal CompressorIn_bh30_160_274 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_160_160 :  std_logic_vector(2 downto 0);
signal heap_bh30_w87_18 :  std_logic;
signal heap_bh30_w88_17 :  std_logic;
signal heap_bh30_w89_15 :  std_logic;
signal CompressorIn_bh30_161_275 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_161_161 :  std_logic_vector(2 downto 0);
signal heap_bh30_w88_18 :  std_logic;
signal heap_bh30_w89_16 :  std_logic;
signal heap_bh30_w90_15 :  std_logic;
signal CompressorIn_bh30_162_276 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_162_162 :  std_logic_vector(2 downto 0);
signal heap_bh30_w89_17 :  std_logic;
signal heap_bh30_w90_16 :  std_logic;
signal heap_bh30_w91_14 :  std_logic;
signal CompressorIn_bh30_163_277 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_163_163 :  std_logic_vector(2 downto 0);
signal heap_bh30_w90_17 :  std_logic;
signal heap_bh30_w91_15 :  std_logic;
signal heap_bh30_w92_11 :  std_logic;
signal CompressorIn_bh30_164_278 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_164_164 :  std_logic_vector(2 downto 0);
signal heap_bh30_w91_16 :  std_logic;
signal heap_bh30_w92_12 :  std_logic;
signal heap_bh30_w93_10 :  std_logic;
signal CompressorIn_bh30_165_279 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_165_165 :  std_logic_vector(2 downto 0);
signal heap_bh30_w92_13 :  std_logic;
signal heap_bh30_w93_11 :  std_logic;
signal heap_bh30_w94_9 :  std_logic;
signal CompressorIn_bh30_166_280 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_166_166 :  std_logic_vector(2 downto 0);
signal heap_bh30_w93_12 :  std_logic;
signal heap_bh30_w94_10 :  std_logic;
signal heap_bh30_w95_8 :  std_logic;
signal CompressorIn_bh30_167_281 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_167_167 :  std_logic_vector(2 downto 0);
signal heap_bh30_w94_11 :  std_logic;
signal heap_bh30_w95_9 :  std_logic;
signal heap_bh30_w96_8 :  std_logic;
signal CompressorIn_bh30_168_282 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_168_168 :  std_logic_vector(2 downto 0);
signal heap_bh30_w95_10 :  std_logic;
signal heap_bh30_w96_9 :  std_logic;
signal heap_bh30_w97_8 :  std_logic;
signal CompressorIn_bh30_169_283 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_169_169 :  std_logic_vector(2 downto 0);
signal heap_bh30_w96_10 :  std_logic;
signal heap_bh30_w97_9 :  std_logic;
signal heap_bh30_w98_8 :  std_logic;
signal CompressorIn_bh30_170_284 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_170_170 :  std_logic_vector(2 downto 0);
signal heap_bh30_w97_10 :  std_logic;
signal heap_bh30_w98_9 :  std_logic;
signal heap_bh30_w99_8 :  std_logic;
signal CompressorIn_bh30_171_285 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_171_171 :  std_logic_vector(2 downto 0);
signal heap_bh30_w98_10 :  std_logic;
signal heap_bh30_w99_9 :  std_logic;
signal heap_bh30_w100_8 :  std_logic;
signal CompressorIn_bh30_172_286 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_172_172 :  std_logic_vector(2 downto 0);
signal heap_bh30_w99_10 :  std_logic;
signal heap_bh30_w100_9 :  std_logic;
signal heap_bh30_w101_8 :  std_logic;
signal CompressorIn_bh30_173_287 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_173_173 :  std_logic_vector(2 downto 0);
signal heap_bh30_w100_10 :  std_logic;
signal heap_bh30_w101_9 :  std_logic;
signal heap_bh30_w102_8 :  std_logic;
signal CompressorIn_bh30_174_288 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_174_174 :  std_logic_vector(2 downto 0);
signal heap_bh30_w101_10 :  std_logic;
signal heap_bh30_w102_9 :  std_logic;
signal heap_bh30_w103_8 :  std_logic;
signal CompressorIn_bh30_175_289 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_175_175 :  std_logic_vector(2 downto 0);
signal heap_bh30_w102_10 :  std_logic;
signal heap_bh30_w103_9 :  std_logic;
signal heap_bh30_w104_8 :  std_logic;
signal CompressorIn_bh30_176_290 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_176_176 :  std_logic_vector(2 downto 0);
signal heap_bh30_w103_10 :  std_logic;
signal heap_bh30_w104_9 :  std_logic;
signal heap_bh30_w105_8 :  std_logic;
signal CompressorIn_bh30_177_291 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_177_177 :  std_logic_vector(2 downto 0);
signal heap_bh30_w104_10 :  std_logic;
signal heap_bh30_w105_9 :  std_logic;
signal heap_bh30_w106_8 :  std_logic;
signal CompressorIn_bh30_178_292 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_178_178 :  std_logic_vector(2 downto 0);
signal heap_bh30_w105_10 :  std_logic;
signal heap_bh30_w106_9 :  std_logic;
signal heap_bh30_w107_8 :  std_logic;
signal CompressorIn_bh30_179_293 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_179_179 :  std_logic_vector(2 downto 0);
signal heap_bh30_w106_10 :  std_logic;
signal heap_bh30_w107_9 :  std_logic;
signal heap_bh30_w108_7 :  std_logic;
signal CompressorIn_bh30_180_294 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_180_180 :  std_logic_vector(2 downto 0);
signal heap_bh30_w107_10 :  std_logic;
signal heap_bh30_w108_8 :  std_logic;
signal heap_bh30_w109_7 :  std_logic;
signal CompressorIn_bh30_181_295 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_181_181 :  std_logic_vector(2 downto 0);
signal heap_bh30_w108_9 :  std_logic;
signal heap_bh30_w109_8 :  std_logic;
signal heap_bh30_w110_7 :  std_logic;
signal CompressorIn_bh30_182_296 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_182_182 :  std_logic_vector(2 downto 0);
signal heap_bh30_w109_9 :  std_logic;
signal heap_bh30_w110_8 :  std_logic;
signal heap_bh30_w111_7 :  std_logic;
signal CompressorIn_bh30_183_297 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_183_183 :  std_logic_vector(2 downto 0);
signal heap_bh30_w110_9 :  std_logic;
signal heap_bh30_w111_8 :  std_logic;
signal heap_bh30_w112_6 :  std_logic;
signal CompressorIn_bh30_184_298 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_184_184 :  std_logic_vector(2 downto 0);
signal heap_bh30_w111_9 :  std_logic;
signal heap_bh30_w112_7 :  std_logic;
signal heap_bh30_w113_6 :  std_logic;
signal CompressorIn_bh30_185_299 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_185_185 :  std_logic_vector(2 downto 0);
signal heap_bh30_w112_8 :  std_logic;
signal heap_bh30_w113_7 :  std_logic;
signal heap_bh30_w114_6 :  std_logic;
signal CompressorIn_bh30_186_300 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_186_186 :  std_logic_vector(2 downto 0);
signal heap_bh30_w113_8 :  std_logic;
signal heap_bh30_w114_7 :  std_logic;
signal heap_bh30_w115_6 :  std_logic;
signal CompressorIn_bh30_187_301 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_187_187 :  std_logic_vector(2 downto 0);
signal heap_bh30_w114_8 :  std_logic;
signal heap_bh30_w115_7 :  std_logic;
signal heap_bh30_w116_6 :  std_logic;
signal CompressorIn_bh30_188_302 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_188_188 :  std_logic_vector(2 downto 0);
signal heap_bh30_w115_8 :  std_logic;
signal heap_bh30_w116_7 :  std_logic;
signal heap_bh30_w117_6 :  std_logic;
signal CompressorIn_bh30_189_303 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_189_189 :  std_logic_vector(2 downto 0);
signal heap_bh30_w116_8 :  std_logic;
signal heap_bh30_w117_7 :  std_logic;
signal heap_bh30_w118_6 :  std_logic;
signal CompressorIn_bh30_190_304 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_190_190 :  std_logic_vector(2 downto 0);
signal heap_bh30_w117_8 :  std_logic;
signal heap_bh30_w118_7 :  std_logic;
signal heap_bh30_w119_6 :  std_logic;
signal CompressorIn_bh30_191_305 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_191_191 :  std_logic_vector(2 downto 0);
signal heap_bh30_w118_8 :  std_logic;
signal heap_bh30_w119_7 :  std_logic;
signal heap_bh30_w120_6 :  std_logic;
signal CompressorIn_bh30_192_306 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_192_192 :  std_logic_vector(2 downto 0);
signal heap_bh30_w119_8 :  std_logic;
signal heap_bh30_w120_7 :  std_logic;
signal heap_bh30_w121_6 :  std_logic;
signal CompressorIn_bh30_193_307 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_193_193 :  std_logic_vector(2 downto 0);
signal heap_bh30_w120_8 :  std_logic;
signal heap_bh30_w121_7 :  std_logic;
signal heap_bh30_w122_6 :  std_logic;
signal CompressorIn_bh30_194_308 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_194_194 :  std_logic_vector(2 downto 0);
signal heap_bh30_w121_8 :  std_logic;
signal heap_bh30_w122_7 :  std_logic;
signal heap_bh30_w123_6 :  std_logic;
signal CompressorIn_bh30_195_309 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_195_195 :  std_logic_vector(2 downto 0);
signal heap_bh30_w122_8 :  std_logic;
signal heap_bh30_w123_7 :  std_logic;
signal heap_bh30_w124_6 :  std_logic;
signal CompressorIn_bh30_196_310 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_196_196 :  std_logic_vector(2 downto 0);
signal heap_bh30_w123_8 :  std_logic;
signal heap_bh30_w124_7 :  std_logic;
signal heap_bh30_w125_6 :  std_logic;
signal CompressorIn_bh30_197_311 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_197_197 :  std_logic_vector(2 downto 0);
signal heap_bh30_w124_8 :  std_logic;
signal heap_bh30_w125_7 :  std_logic;
signal heap_bh30_w126_6 :  std_logic;
signal CompressorIn_bh30_198_312 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_198_198 :  std_logic_vector(2 downto 0);
signal heap_bh30_w125_8 :  std_logic;
signal heap_bh30_w126_7 :  std_logic;
signal heap_bh30_w127_6 :  std_logic;
signal CompressorIn_bh30_199_313 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_199_199 :  std_logic_vector(2 downto 0);
signal heap_bh30_w126_8 :  std_logic;
signal heap_bh30_w127_7 :  std_logic;
signal heap_bh30_w128_6 :  std_logic;
signal CompressorIn_bh30_200_314 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_200_200 :  std_logic_vector(2 downto 0);
signal heap_bh30_w127_8 :  std_logic;
signal heap_bh30_w128_7 :  std_logic;
signal heap_bh30_w129_5 :  std_logic;
signal CompressorIn_bh30_201_315 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_201_201 :  std_logic_vector(2 downto 0);
signal heap_bh30_w128_8 :  std_logic;
signal heap_bh30_w129_6 :  std_logic;
signal heap_bh30_w130_5 :  std_logic;
signal CompressorIn_bh30_202_316 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_202_317 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_202_202 :  std_logic_vector(2 downto 0);
signal heap_bh30_w18_10 :  std_logic;
signal heap_bh30_w19_10 :  std_logic;
signal heap_bh30_w20_9 :  std_logic;
signal CompressorIn_bh30_203_318 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_203_319 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_203_203 :  std_logic_vector(2 downto 0);
signal heap_bh30_w21_10 :  std_logic;
signal heap_bh30_w22_10 :  std_logic;
signal heap_bh30_w23_10 :  std_logic;
signal CompressorIn_bh30_204_320 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_204_321 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_204_204 :  std_logic_vector(2 downto 0);
signal heap_bh30_w23_11 :  std_logic;
signal heap_bh30_w24_11 :  std_logic;
signal heap_bh30_w25_11 :  std_logic;
signal CompressorIn_bh30_205_322 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_205_323 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_205_205 :  std_logic_vector(2 downto 0);
signal heap_bh30_w24_12 :  std_logic;
signal heap_bh30_w25_12 :  std_logic;
signal heap_bh30_w26_10 :  std_logic;
signal CompressorIn_bh30_206_324 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_206_325 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_206_206 :  std_logic_vector(2 downto 0);
signal heap_bh30_w26_11 :  std_logic;
signal heap_bh30_w27_11 :  std_logic;
signal heap_bh30_w28_11 :  std_logic;
signal CompressorIn_bh30_207_326 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_207_327 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_207_207 :  std_logic_vector(2 downto 0);
signal heap_bh30_w27_12 :  std_logic;
signal heap_bh30_w28_12 :  std_logic;
signal heap_bh30_w29_10 :  std_logic;
signal CompressorIn_bh30_208_328 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_208_329 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_208_208 :  std_logic_vector(2 downto 0);
signal heap_bh30_w29_11 :  std_logic;
signal heap_bh30_w30_11 :  std_logic;
signal heap_bh30_w31_11 :  std_logic;
signal CompressorIn_bh30_209_330 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_209_331 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_209_209 :  std_logic_vector(2 downto 0);
signal heap_bh30_w30_12 :  std_logic;
signal heap_bh30_w31_12 :  std_logic;
signal heap_bh30_w32_10 :  std_logic;
signal CompressorIn_bh30_210_332 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_210_333 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_210_210 :  std_logic_vector(2 downto 0);
signal heap_bh30_w34_13 :  std_logic;
signal heap_bh30_w35_12 :  std_logic;
signal heap_bh30_w36_13 :  std_logic;
signal CompressorIn_bh30_211_334 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_211_335 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_211_211 :  std_logic_vector(2 downto 0);
signal heap_bh30_w37_13 :  std_logic;
signal heap_bh30_w38_12 :  std_logic;
signal heap_bh30_w39_13 :  std_logic;
signal CompressorIn_bh30_212_336 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_212_337 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_212_212 :  std_logic_vector(2 downto 0);
signal heap_bh30_w40_13 :  std_logic;
signal heap_bh30_w41_12 :  std_logic;
signal heap_bh30_w42_13 :  std_logic;
signal CompressorIn_bh30_213_338 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_213_339 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_213_213 :  std_logic_vector(2 downto 0);
signal heap_bh30_w43_13 :  std_logic;
signal heap_bh30_w44_12 :  std_logic;
signal heap_bh30_w45_13 :  std_logic;
signal CompressorIn_bh30_214_340 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_214_341 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_214_214 :  std_logic_vector(2 downto 0);
signal heap_bh30_w72_19 :  std_logic;
signal heap_bh30_w73_19 :  std_logic;
signal heap_bh30_w74_18 :  std_logic;
signal CompressorIn_bh30_215_342 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_215_343 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_215_215 :  std_logic_vector(2 downto 0);
signal heap_bh30_w75_19 :  std_logic;
signal heap_bh30_w76_19 :  std_logic;
signal heap_bh30_w77_18 :  std_logic;
signal CompressorIn_bh30_216_344 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_216_345 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_216_216 :  std_logic_vector(2 downto 0);
signal heap_bh30_w78_19 :  std_logic;
signal heap_bh30_w79_19 :  std_logic;
signal heap_bh30_w80_18 :  std_logic;
signal CompressorIn_bh30_217_346 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_217_347 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_217_217 :  std_logic_vector(2 downto 0);
signal heap_bh30_w81_19 :  std_logic;
signal heap_bh30_w82_19 :  std_logic;
signal heap_bh30_w83_18 :  std_logic;
signal CompressorIn_bh30_218_348 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_218_349 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_218_218 :  std_logic_vector(2 downto 0);
signal heap_bh30_w84_19 :  std_logic;
signal heap_bh30_w85_19 :  std_logic;
signal heap_bh30_w86_18 :  std_logic;
signal CompressorIn_bh30_219_350 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_219_351 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_219_219 :  std_logic_vector(2 downto 0);
signal heap_bh30_w87_19 :  std_logic;
signal heap_bh30_w88_19 :  std_logic;
signal heap_bh30_w89_18 :  std_logic;
signal CompressorIn_bh30_220_352 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_220_353 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_220_220 :  std_logic_vector(2 downto 0);
signal heap_bh30_w90_18 :  std_logic;
signal heap_bh30_w91_17 :  std_logic;
signal heap_bh30_w92_14 :  std_logic;
signal CompressorIn_bh30_221_354 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_221_355 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_221_221 :  std_logic_vector(2 downto 0);
signal heap_bh30_w93_13 :  std_logic;
signal heap_bh30_w94_12 :  std_logic;
signal heap_bh30_w95_11 :  std_logic;
signal CompressorIn_bh30_222_356 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_222_357 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_222_222 :  std_logic_vector(2 downto 0);
signal heap_bh30_w129_7 :  std_logic;
signal heap_bh30_w130_6 :  std_logic;
signal heap_bh30_w131_5 :  std_logic;
signal CompressorIn_bh30_223_358 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_223_359 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_223_223 :  std_logic_vector(2 downto 0);
signal heap_bh30_w130_7 :  std_logic;
signal heap_bh30_w131_6 :  std_logic;
signal heap_bh30_w132_4 :  std_logic;
signal CompressorIn_bh30_224_360 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_224_361 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_224_224 :  std_logic_vector(2 downto 0);
signal heap_bh30_w131_7 :  std_logic;
signal heap_bh30_w132_5 :  std_logic;
signal heap_bh30_w133_4 :  std_logic;
signal CompressorIn_bh30_225_362 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_225_363 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_225_225 :  std_logic_vector(2 downto 0);
signal heap_bh30_w133_5 :  std_logic;
signal heap_bh30_w134_4 :  std_logic;
signal heap_bh30_w135_4 :  std_logic;
signal CompressorIn_bh30_226_364 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_226_365 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_226_226 :  std_logic_vector(2 downto 0);
signal heap_bh30_w135_5 :  std_logic;
signal heap_bh30_w136_4 :  std_logic;
signal heap_bh30_w137_4 :  std_logic;
signal CompressorIn_bh30_227_366 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_227_367 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_227_227 :  std_logic_vector(2 downto 0);
signal heap_bh30_w137_5 :  std_logic;
signal heap_bh30_w138_4 :  std_logic;
signal heap_bh30_w139_4 :  std_logic;
signal CompressorIn_bh30_228_368 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_228_369 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_228_228 :  std_logic_vector(2 downto 0);
signal heap_bh30_w139_5 :  std_logic;
signal heap_bh30_w140_4 :  std_logic;
signal heap_bh30_w141_4 :  std_logic;
signal CompressorIn_bh30_229_370 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_229_371 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_229_229 :  std_logic_vector(2 downto 0);
signal heap_bh30_w141_5 :  std_logic;
signal heap_bh30_w142_4 :  std_logic;
signal heap_bh30_w143_4 :  std_logic;
signal CompressorIn_bh30_230_372 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_230_373 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_230_230 :  std_logic_vector(2 downto 0);
signal heap_bh30_w143_5 :  std_logic;
signal heap_bh30_w144_4 :  std_logic;
signal heap_bh30_w145_4 :  std_logic;
signal CompressorIn_bh30_231_374 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_231_375 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_231_231 :  std_logic_vector(2 downto 0);
signal heap_bh30_w145_5 :  std_logic;
signal heap_bh30_w146_3 :  std_logic;
signal heap_bh30_w147_3 :  std_logic;
signal CompressorIn_bh30_232_376 :  std_logic_vector(4 downto 0);
signal CompressorOut_bh30_232_232 :  std_logic_vector(2 downto 0);
signal heap_bh30_w46_13 :  std_logic;
signal heap_bh30_w47_14 :  std_logic;
signal heap_bh30_w48_15 :  std_logic;
signal CompressorIn_bh30_233_377 :  std_logic_vector(3 downto 0);
signal CompressorOut_bh30_233_233 :  std_logic_vector(2 downto 0);
signal heap_bh30_w32_11 :  std_logic;
signal heap_bh30_w33_13 :  std_logic;
signal heap_bh30_w34_14 :  std_logic;
signal CompressorIn_bh30_234_378 :  std_logic_vector(3 downto 0);
signal CompressorOut_bh30_234_234 :  std_logic_vector(2 downto 0);
signal heap_bh30_w35_13 :  std_logic;
signal heap_bh30_w36_14 :  std_logic;
signal heap_bh30_w37_14 :  std_logic;
signal CompressorIn_bh30_235_379 :  std_logic_vector(3 downto 0);
signal CompressorOut_bh30_235_235 :  std_logic_vector(2 downto 0);
signal heap_bh30_w38_13 :  std_logic;
signal heap_bh30_w39_14 :  std_logic;
signal heap_bh30_w40_14 :  std_logic;
signal CompressorIn_bh30_236_380 :  std_logic_vector(3 downto 0);
signal CompressorOut_bh30_236_236 :  std_logic_vector(2 downto 0);
signal heap_bh30_w41_13 :  std_logic;
signal heap_bh30_w42_14 :  std_logic;
signal heap_bh30_w43_14 :  std_logic;
signal CompressorIn_bh30_237_381 :  std_logic_vector(3 downto 0);
signal CompressorOut_bh30_237_237 :  std_logic_vector(2 downto 0);
signal heap_bh30_w44_13 :  std_logic;
signal heap_bh30_w45_14 :  std_logic;
signal heap_bh30_w46_14 :  std_logic;
signal CompressorIn_bh30_238_382 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_238_383 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_238_238 :  std_logic_vector(2 downto 0);
signal heap_bh30_w2_3 :  std_logic;
signal heap_bh30_w3_5 :  std_logic;
signal heap_bh30_w4_5 :  std_logic;
signal CompressorIn_bh30_239_384 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_239_385 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_239_239 :  std_logic_vector(2 downto 0);
signal heap_bh30_w4_6 :  std_logic;
signal heap_bh30_w5_6 :  std_logic;
signal heap_bh30_w6_7 :  std_logic;
signal CompressorIn_bh30_240_386 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_240_387 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_240_240 :  std_logic_vector(2 downto 0);
signal heap_bh30_w6_8 :  std_logic;
signal heap_bh30_w7_7 :  std_logic;
signal heap_bh30_w8_7 :  std_logic;
signal CompressorIn_bh30_241_388 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_241_389 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_241_241 :  std_logic_vector(2 downto 0);
signal heap_bh30_w12_9 :  std_logic;
signal heap_bh30_w13_9 :  std_logic;
signal heap_bh30_w14_8 :  std_logic;
signal CompressorIn_bh30_242_390 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_242_391 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_242_242 :  std_logic_vector(2 downto 0);
signal heap_bh30_w15_9 :  std_logic;
signal heap_bh30_w16_10 :  std_logic;
signal heap_bh30_w17_9 :  std_logic;
signal CompressorIn_bh30_243_392 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_243_393 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_243_243 :  std_logic_vector(2 downto 0);
signal heap_bh30_w69_18 :  std_logic;
signal heap_bh30_w70_18 :  std_logic;
signal heap_bh30_w71_18 :  std_logic;
signal CompressorIn_bh30_244_394 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_244_395 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_244_244 :  std_logic_vector(2 downto 0);
signal heap_bh30_w147_4 :  std_logic;
signal heap_bh30_w148_3 :  std_logic;
signal heap_bh30_w149_3 :  std_logic;
signal CompressorIn_bh30_245_396 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_245_397 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_245_245 :  std_logic_vector(2 downto 0);
signal heap_bh30_w149_4 :  std_logic;
signal heap_bh30_w150_3 :  std_logic;
signal heap_bh30_w151_3 :  std_logic;
signal CompressorIn_bh30_246_398 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_246_399 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_246_246 :  std_logic_vector(2 downto 0);
signal heap_bh30_w151_4 :  std_logic;
signal heap_bh30_w152_3 :  std_logic;
signal heap_bh30_w153_3 :  std_logic;
signal CompressorIn_bh30_247_400 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_247_401 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_247_247 :  std_logic_vector(2 downto 0);
signal heap_bh30_w153_4 :  std_logic;
signal heap_bh30_w154_3 :  std_logic;
signal heap_bh30_w155_3 :  std_logic;
signal CompressorIn_bh30_248_402 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_248_403 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_248_248 :  std_logic_vector(2 downto 0);
signal heap_bh30_w155_4 :  std_logic;
signal heap_bh30_w156_2 :  std_logic;
signal heap_bh30_w157_2 :  std_logic;
signal CompressorIn_bh30_249_404 :  std_logic_vector(2 downto 0);
signal CompressorOut_bh30_249_249 :  std_logic_vector(1 downto 0);
signal heap_bh30_w17_10 :  std_logic;
signal heap_bh30_w18_11 :  std_logic;
signal CompressorIn_bh30_250_405 :  std_logic_vector(2 downto 0);
signal CompressorOut_bh30_250_250 :  std_logic_vector(1 downto 0);
signal heap_bh30_w20_10 :  std_logic;
signal heap_bh30_w21_11 :  std_logic;
signal CompressorIn_bh30_251_406 :  std_logic_vector(2 downto 0);
signal CompressorOut_bh30_251_251 :  std_logic_vector(1 downto 0);
signal heap_bh30_w25_13 :  std_logic;
signal heap_bh30_w26_12 :  std_logic;
signal CompressorIn_bh30_252_407 :  std_logic_vector(2 downto 0);
signal CompressorOut_bh30_252_252 :  std_logic_vector(1 downto 0);
signal heap_bh30_w28_13 :  std_logic;
signal heap_bh30_w29_12 :  std_logic;
signal CompressorIn_bh30_253_408 :  std_logic_vector(2 downto 0);
signal CompressorOut_bh30_253_253 :  std_logic_vector(1 downto 0);
signal heap_bh30_w31_13 :  std_logic;
signal heap_bh30_w32_12 :  std_logic;
signal CompressorIn_bh30_254_409 :  std_logic_vector(2 downto 0);
signal CompressorOut_bh30_254_254 :  std_logic_vector(1 downto 0);
signal heap_bh30_w71_19 :  std_logic;
signal heap_bh30_w72_20 :  std_logic;
signal CompressorIn_bh30_255_410 :  std_logic_vector(2 downto 0);
signal CompressorOut_bh30_255_255 :  std_logic_vector(1 downto 0);
signal heap_bh30_w74_19 :  std_logic;
signal heap_bh30_w75_20 :  std_logic;
signal CompressorIn_bh30_256_411 :  std_logic_vector(2 downto 0);
signal CompressorOut_bh30_256_256 :  std_logic_vector(1 downto 0);
signal heap_bh30_w77_19 :  std_logic;
signal heap_bh30_w78_20 :  std_logic;
signal CompressorIn_bh30_257_412 :  std_logic_vector(2 downto 0);
signal CompressorOut_bh30_257_257 :  std_logic_vector(1 downto 0);
signal heap_bh30_w80_19 :  std_logic;
signal heap_bh30_w81_20 :  std_logic;
signal CompressorIn_bh30_258_413 :  std_logic_vector(2 downto 0);
signal CompressorOut_bh30_258_258 :  std_logic_vector(1 downto 0);
signal heap_bh30_w83_19 :  std_logic;
signal heap_bh30_w84_20 :  std_logic;
signal CompressorIn_bh30_259_414 :  std_logic_vector(2 downto 0);
signal CompressorOut_bh30_259_259 :  std_logic_vector(1 downto 0);
signal heap_bh30_w86_19 :  std_logic;
signal heap_bh30_w87_20 :  std_logic;
signal CompressorIn_bh30_260_415 :  std_logic_vector(2 downto 0);
signal CompressorOut_bh30_260_260 :  std_logic_vector(1 downto 0);
signal heap_bh30_w89_19 :  std_logic;
signal heap_bh30_w90_19 :  std_logic;
signal CompressorIn_bh30_261_416 :  std_logic_vector(2 downto 0);
signal CompressorOut_bh30_261_261 :  std_logic_vector(1 downto 0);
signal heap_bh30_w92_15 :  std_logic;
signal heap_bh30_w93_14 :  std_logic;
signal CompressorIn_bh30_262_417 :  std_logic_vector(2 downto 0);
signal CompressorOut_bh30_262_262 :  std_logic_vector(1 downto 0);
signal heap_bh30_w132_6 :  std_logic;
signal heap_bh30_w133_6 :  std_logic;
signal CompressorIn_bh30_263_418 :  std_logic_vector(2 downto 0);
signal CompressorOut_bh30_263_263 :  std_logic_vector(1 downto 0);
signal heap_bh30_w134_5 :  std_logic;
signal heap_bh30_w135_6 :  std_logic;
signal CompressorIn_bh30_264_419 :  std_logic_vector(2 downto 0);
signal CompressorOut_bh30_264_264 :  std_logic_vector(1 downto 0);
signal heap_bh30_w136_5 :  std_logic;
signal heap_bh30_w137_6 :  std_logic;
signal CompressorIn_bh30_265_420 :  std_logic_vector(2 downto 0);
signal CompressorOut_bh30_265_265 :  std_logic_vector(1 downto 0);
signal heap_bh30_w138_5 :  std_logic;
signal heap_bh30_w139_6 :  std_logic;
signal CompressorIn_bh30_266_421 :  std_logic_vector(2 downto 0);
signal CompressorOut_bh30_266_266 :  std_logic_vector(1 downto 0);
signal heap_bh30_w140_5 :  std_logic;
signal heap_bh30_w141_6 :  std_logic;
signal CompressorIn_bh30_267_422 :  std_logic_vector(2 downto 0);
signal CompressorOut_bh30_267_267 :  std_logic_vector(1 downto 0);
signal heap_bh30_w142_5 :  std_logic;
signal heap_bh30_w143_6 :  std_logic;
signal CompressorIn_bh30_268_423 :  std_logic_vector(2 downto 0);
signal CompressorOut_bh30_268_268 :  std_logic_vector(1 downto 0);
signal heap_bh30_w144_5 :  std_logic;
signal heap_bh30_w145_6 :  std_logic;
signal CompressorIn_bh30_269_424 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_269_269 :  std_logic_vector(2 downto 0);
signal heap_bh30_w73_20 :  std_logic;
signal heap_bh30_w74_20 :  std_logic;
signal heap_bh30_w75_21 :  std_logic;
signal CompressorIn_bh30_270_425 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_270_270 :  std_logic_vector(2 downto 0);
signal heap_bh30_w76_20 :  std_logic;
signal heap_bh30_w77_20 :  std_logic;
signal heap_bh30_w78_21 :  std_logic;
signal CompressorIn_bh30_271_426 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_271_271 :  std_logic_vector(2 downto 0);
signal heap_bh30_w79_20 :  std_logic;
signal heap_bh30_w80_20 :  std_logic;
signal heap_bh30_w81_21 :  std_logic;
signal CompressorIn_bh30_272_427 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_272_272 :  std_logic_vector(2 downto 0);
signal heap_bh30_w82_20 :  std_logic;
signal heap_bh30_w83_20 :  std_logic;
signal heap_bh30_w84_21 :  std_logic;
signal CompressorIn_bh30_273_428 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_273_273 :  std_logic_vector(2 downto 0);
signal heap_bh30_w85_20 :  std_logic;
signal heap_bh30_w86_20 :  std_logic;
signal heap_bh30_w87_21 :  std_logic;
signal CompressorIn_bh30_274_429 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_274_274 :  std_logic_vector(2 downto 0);
signal heap_bh30_w88_20 :  std_logic;
signal heap_bh30_w89_20 :  std_logic;
signal heap_bh30_w90_20 :  std_logic;
signal CompressorIn_bh30_275_430 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_275_275 :  std_logic_vector(2 downto 0);
signal heap_bh30_w91_18 :  std_logic;
signal heap_bh30_w92_16 :  std_logic;
signal heap_bh30_w93_15 :  std_logic;
signal CompressorIn_bh30_276_431 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_276_276 :  std_logic_vector(2 downto 0);
signal heap_bh30_w94_13 :  std_logic;
signal heap_bh30_w95_12 :  std_logic;
signal heap_bh30_w96_11 :  std_logic;
signal CompressorIn_bh30_277_432 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_277_277 :  std_logic_vector(2 downto 0);
signal heap_bh30_w95_13 :  std_logic;
signal heap_bh30_w96_12 :  std_logic;
signal heap_bh30_w97_11 :  std_logic;
signal CompressorIn_bh30_278_433 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_278_434 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_278_278 :  std_logic_vector(2 downto 0);
signal heap_bh30_w34_15 :  std_logic;
signal heap_bh30_w35_14 :  std_logic;
signal heap_bh30_w36_15 :  std_logic;
signal CompressorIn_bh30_279_435 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_279_436 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_279_279 :  std_logic_vector(2 downto 0);
signal heap_bh30_w37_15 :  std_logic;
signal heap_bh30_w38_14 :  std_logic;
signal heap_bh30_w39_15 :  std_logic;
signal CompressorIn_bh30_280_437 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_280_438 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_280_280 :  std_logic_vector(2 downto 0);
signal heap_bh30_w40_15 :  std_logic;
signal heap_bh30_w41_14 :  std_logic;
signal heap_bh30_w42_15 :  std_logic;
signal CompressorIn_bh30_281_439 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_281_440 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_281_281 :  std_logic_vector(2 downto 0);
signal heap_bh30_w43_15 :  std_logic;
signal heap_bh30_w44_14 :  std_logic;
signal heap_bh30_w45_15 :  std_logic;
signal CompressorIn_bh30_282_441 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_282_442 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_282_282 :  std_logic_vector(2 downto 0);
signal heap_bh30_w48_16 :  std_logic;
signal heap_bh30_w49_16 :  std_logic;
signal heap_bh30_w50_16 :  std_logic;
signal CompressorIn_bh30_283_443 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_283_444 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_283_283 :  std_logic_vector(2 downto 0);
signal heap_bh30_w50_17 :  std_logic;
signal heap_bh30_w51_17 :  std_logic;
signal heap_bh30_w52_17 :  std_logic;
signal CompressorIn_bh30_284_445 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_284_446 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_284_284 :  std_logic_vector(2 downto 0);
signal heap_bh30_w51_18 :  std_logic;
signal heap_bh30_w52_18 :  std_logic;
signal heap_bh30_w53_16 :  std_logic;
signal CompressorIn_bh30_285_447 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_285_448 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_285_285 :  std_logic_vector(2 downto 0);
signal heap_bh30_w53_17 :  std_logic;
signal heap_bh30_w54_17 :  std_logic;
signal heap_bh30_w55_17 :  std_logic;
signal CompressorIn_bh30_286_449 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_286_450 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_286_286 :  std_logic_vector(2 downto 0);
signal heap_bh30_w54_18 :  std_logic;
signal heap_bh30_w55_18 :  std_logic;
signal heap_bh30_w56_16 :  std_logic;
signal CompressorIn_bh30_287_451 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_287_452 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_287_287 :  std_logic_vector(2 downto 0);
signal heap_bh30_w56_17 :  std_logic;
signal heap_bh30_w57_17 :  std_logic;
signal heap_bh30_w58_17 :  std_logic;
signal CompressorIn_bh30_288_453 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_288_454 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_288_288 :  std_logic_vector(2 downto 0);
signal heap_bh30_w57_18 :  std_logic;
signal heap_bh30_w58_18 :  std_logic;
signal heap_bh30_w59_16 :  std_logic;
signal CompressorIn_bh30_289_455 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_289_456 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_289_289 :  std_logic_vector(2 downto 0);
signal heap_bh30_w59_17 :  std_logic;
signal heap_bh30_w60_17 :  std_logic;
signal heap_bh30_w61_17 :  std_logic;
signal CompressorIn_bh30_290_457 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_290_458 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_290_290 :  std_logic_vector(2 downto 0);
signal heap_bh30_w60_18 :  std_logic;
signal heap_bh30_w61_18 :  std_logic;
signal heap_bh30_w62_16 :  std_logic;
signal CompressorIn_bh30_291_459 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_291_460 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_291_291 :  std_logic_vector(2 downto 0);
signal heap_bh30_w62_17 :  std_logic;
signal heap_bh30_w63_17 :  std_logic;
signal heap_bh30_w64_17 :  std_logic;
signal CompressorIn_bh30_292_461 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_292_462 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_292_292 :  std_logic_vector(2 downto 0);
signal heap_bh30_w63_18 :  std_logic;
signal heap_bh30_w64_18 :  std_logic;
signal heap_bh30_w65_16 :  std_logic;
signal CompressorIn_bh30_293_463 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_293_464 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_293_293 :  std_logic_vector(2 downto 0);
signal heap_bh30_w65_17 :  std_logic;
signal heap_bh30_w66_17 :  std_logic;
signal heap_bh30_w67_18 :  std_logic;
signal CompressorIn_bh30_294_465 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_294_466 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_294_294 :  std_logic_vector(2 downto 0);
signal heap_bh30_w66_18 :  std_logic;
signal heap_bh30_w67_19 :  std_logic;
signal heap_bh30_w68_17 :  std_logic;
signal CompressorIn_bh30_295_467 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_295_468 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_295_295 :  std_logic_vector(2 downto 0);
signal heap_bh30_w67_20 :  std_logic;
signal heap_bh30_w68_18 :  std_logic;
signal heap_bh30_w69_19 :  std_logic;
signal CompressorIn_bh30_296_469 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_296_470 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_296_296 :  std_logic_vector(2 downto 0);
signal heap_bh30_w68_19 :  std_logic;
signal heap_bh30_w69_20 :  std_logic;
signal heap_bh30_w70_19 :  std_logic;
signal CompressorIn_bh30_297_471 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_297_472 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_297_297 :  std_logic_vector(2 downto 0);
signal heap_bh30_w70_20 :  std_logic;
signal heap_bh30_w71_20 :  std_logic;
signal heap_bh30_w72_21 :  std_logic;
signal CompressorIn_bh30_298_473 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_298_474 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_298_298 :  std_logic_vector(2 downto 0);
signal heap_bh30_w71_21 :  std_logic;
signal heap_bh30_w72_22 :  std_logic;
signal heap_bh30_w73_21 :  std_logic;
signal CompressorIn_bh30_299_475 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_299_476 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_299_299 :  std_logic_vector(2 downto 0);
signal heap_bh30_w74_21 :  std_logic;
signal heap_bh30_w75_22 :  std_logic;
signal heap_bh30_w76_21 :  std_logic;
signal CompressorIn_bh30_300_477 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_300_478 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_300_300 :  std_logic_vector(2 downto 0);
signal heap_bh30_w77_21 :  std_logic;
signal heap_bh30_w78_22 :  std_logic;
signal heap_bh30_w79_21 :  std_logic;
signal CompressorIn_bh30_301_479 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_301_480 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_301_301 :  std_logic_vector(2 downto 0);
signal heap_bh30_w80_21 :  std_logic;
signal heap_bh30_w81_22 :  std_logic;
signal heap_bh30_w82_21 :  std_logic;
signal CompressorIn_bh30_302_481 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_302_482 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_302_302 :  std_logic_vector(2 downto 0);
signal heap_bh30_w83_21 :  std_logic;
signal heap_bh30_w84_22 :  std_logic;
signal heap_bh30_w85_21 :  std_logic;
signal CompressorIn_bh30_303_483 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_303_484 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_303_303 :  std_logic_vector(2 downto 0);
signal heap_bh30_w86_21 :  std_logic;
signal heap_bh30_w87_22 :  std_logic;
signal heap_bh30_w88_21 :  std_logic;
signal CompressorIn_bh30_304_485 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_304_486 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_304_304 :  std_logic_vector(2 downto 0);
signal heap_bh30_w89_21 :  std_logic;
signal heap_bh30_w90_21 :  std_logic;
signal heap_bh30_w91_19 :  std_logic;
signal CompressorIn_bh30_305_487 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_305_488 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_305_305 :  std_logic_vector(2 downto 0);
signal heap_bh30_w92_17 :  std_logic;
signal heap_bh30_w93_16 :  std_logic;
signal heap_bh30_w94_14 :  std_logic;
signal CompressorIn_bh30_306_489 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_306_490 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_306_306 :  std_logic_vector(2 downto 0);
signal heap_bh30_w96_13 :  std_logic;
signal heap_bh30_w97_12 :  std_logic;
signal heap_bh30_w98_11 :  std_logic;
signal CompressorIn_bh30_307_491 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_307_492 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_307_307 :  std_logic_vector(2 downto 0);
signal heap_bh30_w97_13 :  std_logic;
signal heap_bh30_w98_12 :  std_logic;
signal heap_bh30_w99_11 :  std_logic;
signal CompressorIn_bh30_308_493 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_308_494 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_308_308 :  std_logic_vector(2 downto 0);
signal heap_bh30_w98_13 :  std_logic;
signal heap_bh30_w99_12 :  std_logic;
signal heap_bh30_w100_11 :  std_logic;
signal CompressorIn_bh30_309_495 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_309_496 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_309_309 :  std_logic_vector(2 downto 0);
signal heap_bh30_w99_13 :  std_logic;
signal heap_bh30_w100_12 :  std_logic;
signal heap_bh30_w101_11 :  std_logic;
signal CompressorIn_bh30_310_497 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_310_498 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_310_310 :  std_logic_vector(2 downto 0);
signal heap_bh30_w100_13 :  std_logic;
signal heap_bh30_w101_12 :  std_logic;
signal heap_bh30_w102_11 :  std_logic;
signal CompressorIn_bh30_311_499 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_311_500 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_311_311 :  std_logic_vector(2 downto 0);
signal heap_bh30_w101_13 :  std_logic;
signal heap_bh30_w102_12 :  std_logic;
signal heap_bh30_w103_11 :  std_logic;
signal CompressorIn_bh30_312_501 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_312_502 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_312_312 :  std_logic_vector(2 downto 0);
signal heap_bh30_w102_13 :  std_logic;
signal heap_bh30_w103_12 :  std_logic;
signal heap_bh30_w104_11 :  std_logic;
signal CompressorIn_bh30_313_503 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_313_504 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_313_313 :  std_logic_vector(2 downto 0);
signal heap_bh30_w103_13 :  std_logic;
signal heap_bh30_w104_12 :  std_logic;
signal heap_bh30_w105_11 :  std_logic;
signal CompressorIn_bh30_314_505 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_314_506 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_314_314 :  std_logic_vector(2 downto 0);
signal heap_bh30_w104_13 :  std_logic;
signal heap_bh30_w105_12 :  std_logic;
signal heap_bh30_w106_11 :  std_logic;
signal CompressorIn_bh30_315_507 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_315_508 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_315_315 :  std_logic_vector(2 downto 0);
signal heap_bh30_w105_13 :  std_logic;
signal heap_bh30_w106_12 :  std_logic;
signal heap_bh30_w107_11 :  std_logic;
signal CompressorIn_bh30_316_509 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_316_510 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_316_316 :  std_logic_vector(2 downto 0);
signal heap_bh30_w106_13 :  std_logic;
signal heap_bh30_w107_12 :  std_logic;
signal heap_bh30_w108_10 :  std_logic;
signal CompressorIn_bh30_317_511 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_317_512 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_317_317 :  std_logic_vector(2 downto 0);
signal heap_bh30_w107_13 :  std_logic;
signal heap_bh30_w108_11 :  std_logic;
signal heap_bh30_w109_10 :  std_logic;
signal CompressorIn_bh30_318_513 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_318_514 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_318_318 :  std_logic_vector(2 downto 0);
signal heap_bh30_w109_11 :  std_logic;
signal heap_bh30_w110_10 :  std_logic;
signal heap_bh30_w111_10 :  std_logic;
signal CompressorIn_bh30_319_515 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_319_516 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_319_319 :  std_logic_vector(2 downto 0);
signal heap_bh30_w111_11 :  std_logic;
signal heap_bh30_w112_9 :  std_logic;
signal heap_bh30_w113_9 :  std_logic;
signal CompressorIn_bh30_320_517 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_320_518 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_320_320 :  std_logic_vector(2 downto 0);
signal heap_bh30_w129_8 :  std_logic;
signal heap_bh30_w130_8 :  std_logic;
signal heap_bh30_w131_8 :  std_logic;
signal CompressorIn_bh30_321_519 :  std_logic_vector(3 downto 0);
signal CompressorOut_bh30_321_321 :  std_logic_vector(2 downto 0);
signal heap_bh30_w72_23 :  std_logic;
signal heap_bh30_w73_22 :  std_logic;
signal heap_bh30_w74_22 :  std_logic;
signal CompressorIn_bh30_322_520 :  std_logic_vector(3 downto 0);
signal CompressorOut_bh30_322_322 :  std_logic_vector(2 downto 0);
signal heap_bh30_w75_23 :  std_logic;
signal heap_bh30_w76_22 :  std_logic;
signal heap_bh30_w77_22 :  std_logic;
signal CompressorIn_bh30_323_521 :  std_logic_vector(3 downto 0);
signal CompressorOut_bh30_323_323 :  std_logic_vector(2 downto 0);
signal heap_bh30_w78_23 :  std_logic;
signal heap_bh30_w79_22 :  std_logic;
signal heap_bh30_w80_22 :  std_logic;
signal CompressorIn_bh30_324_522 :  std_logic_vector(3 downto 0);
signal CompressorOut_bh30_324_324 :  std_logic_vector(2 downto 0);
signal heap_bh30_w81_23 :  std_logic;
signal heap_bh30_w82_22 :  std_logic;
signal heap_bh30_w83_22 :  std_logic;
signal CompressorIn_bh30_325_523 :  std_logic_vector(3 downto 0);
signal CompressorOut_bh30_325_325 :  std_logic_vector(2 downto 0);
signal heap_bh30_w84_23 :  std_logic;
signal heap_bh30_w85_22 :  std_logic;
signal heap_bh30_w86_22 :  std_logic;
signal CompressorIn_bh30_326_524 :  std_logic_vector(3 downto 0);
signal CompressorOut_bh30_326_326 :  std_logic_vector(2 downto 0);
signal heap_bh30_w87_23 :  std_logic;
signal heap_bh30_w88_22 :  std_logic;
signal heap_bh30_w89_22 :  std_logic;
signal CompressorIn_bh30_327_525 :  std_logic_vector(3 downto 0);
signal CompressorOut_bh30_327_327 :  std_logic_vector(2 downto 0);
signal heap_bh30_w90_22 :  std_logic;
signal heap_bh30_w91_20 :  std_logic;
signal heap_bh30_w92_18 :  std_logic;
signal CompressorIn_bh30_328_526 :  std_logic_vector(3 downto 0);
signal CompressorOut_bh30_328_328 :  std_logic_vector(2 downto 0);
signal heap_bh30_w93_17 :  std_logic;
signal heap_bh30_w94_15 :  std_logic;
signal heap_bh30_w95_14 :  std_logic;
signal CompressorIn_bh30_329_527 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_329_528 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_329_329 :  std_logic_vector(2 downto 0);
signal heap_bh30_w8_8 :  std_logic;
signal heap_bh30_w9_8 :  std_logic;
signal heap_bh30_w10_9 :  std_logic;
signal CompressorIn_bh30_330_529 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_330_530 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_330_330 :  std_logic_vector(2 downto 0);
signal heap_bh30_w19_11 :  std_logic;
signal heap_bh30_w20_11 :  std_logic;
signal heap_bh30_w21_12 :  std_logic;
signal CompressorIn_bh30_331_531 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_331_532 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_331_331 :  std_logic_vector(2 downto 0);
signal heap_bh30_w22_11 :  std_logic;
signal heap_bh30_w23_12 :  std_logic;
signal heap_bh30_w24_13 :  std_logic;
signal CompressorIn_bh30_332_533 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_332_534 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_332_332 :  std_logic_vector(2 downto 0);
signal heap_bh30_w25_14 :  std_logic;
signal heap_bh30_w26_13 :  std_logic;
signal heap_bh30_w27_13 :  std_logic;
signal CompressorIn_bh30_333_535 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_333_536 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_333_333 :  std_logic_vector(2 downto 0);
signal heap_bh30_w28_14 :  std_logic;
signal heap_bh30_w29_13 :  std_logic;
signal heap_bh30_w30_13 :  std_logic;
signal CompressorIn_bh30_334_537 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_334_538 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_334_334 :  std_logic_vector(2 downto 0);
signal heap_bh30_w31_14 :  std_logic;
signal heap_bh30_w32_13 :  std_logic;
signal heap_bh30_w33_14 :  std_logic;
signal CompressorIn_bh30_335_539 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_335_540 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_335_335 :  std_logic_vector(2 downto 0);
signal heap_bh30_w45_16 :  std_logic;
signal heap_bh30_w46_15 :  std_logic;
signal heap_bh30_w47_15 :  std_logic;
signal CompressorIn_bh30_336_541 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_336_542 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_336_336 :  std_logic_vector(2 downto 0);
signal heap_bh30_w113_10 :  std_logic;
signal heap_bh30_w114_9 :  std_logic;
signal heap_bh30_w115_9 :  std_logic;
signal CompressorIn_bh30_337_543 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_337_544 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_337_337 :  std_logic_vector(2 downto 0);
signal heap_bh30_w115_10 :  std_logic;
signal heap_bh30_w116_9 :  std_logic;
signal heap_bh30_w117_9 :  std_logic;
signal CompressorIn_bh30_338_545 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_338_546 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_338_338 :  std_logic_vector(2 downto 0);
signal heap_bh30_w117_10 :  std_logic;
signal heap_bh30_w118_9 :  std_logic;
signal heap_bh30_w119_9 :  std_logic;
signal CompressorIn_bh30_339_547 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_339_548 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_339_339 :  std_logic_vector(2 downto 0);
signal heap_bh30_w119_10 :  std_logic;
signal heap_bh30_w120_9 :  std_logic;
signal heap_bh30_w121_9 :  std_logic;
signal CompressorIn_bh30_340_549 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_340_550 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_340_340 :  std_logic_vector(2 downto 0);
signal heap_bh30_w121_10 :  std_logic;
signal heap_bh30_w122_9 :  std_logic;
signal heap_bh30_w123_9 :  std_logic;
signal CompressorIn_bh30_341_551 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_341_552 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_341_341 :  std_logic_vector(2 downto 0);
signal heap_bh30_w123_10 :  std_logic;
signal heap_bh30_w124_9 :  std_logic;
signal heap_bh30_w125_9 :  std_logic;
signal CompressorIn_bh30_342_553 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_342_554 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_342_342 :  std_logic_vector(2 downto 0);
signal heap_bh30_w125_10 :  std_logic;
signal heap_bh30_w126_9 :  std_logic;
signal heap_bh30_w127_9 :  std_logic;
signal CompressorIn_bh30_343_555 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_343_556 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_343_343 :  std_logic_vector(2 downto 0);
signal heap_bh30_w127_10 :  std_logic;
signal heap_bh30_w128_9 :  std_logic;
signal heap_bh30_w129_9 :  std_logic;
signal CompressorIn_bh30_344_557 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_344_558 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_344_344 :  std_logic_vector(2 downto 0);
signal heap_bh30_w131_9 :  std_logic;
signal heap_bh30_w132_7 :  std_logic;
signal heap_bh30_w133_7 :  std_logic;
signal CompressorIn_bh30_345_559 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_345_560 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_345_345 :  std_logic_vector(2 downto 0);
signal heap_bh30_w133_8 :  std_logic;
signal heap_bh30_w134_6 :  std_logic;
signal heap_bh30_w135_7 :  std_logic;
signal CompressorIn_bh30_346_561 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_346_562 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_346_346 :  std_logic_vector(2 downto 0);
signal heap_bh30_w135_8 :  std_logic;
signal heap_bh30_w136_6 :  std_logic;
signal heap_bh30_w137_7 :  std_logic;
signal CompressorIn_bh30_347_563 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_347_564 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_347_347 :  std_logic_vector(2 downto 0);
signal heap_bh30_w137_8 :  std_logic;
signal heap_bh30_w138_6 :  std_logic;
signal heap_bh30_w139_7 :  std_logic;
signal CompressorIn_bh30_348_565 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_348_566 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_348_348 :  std_logic_vector(2 downto 0);
signal heap_bh30_w139_8 :  std_logic;
signal heap_bh30_w140_6 :  std_logic;
signal heap_bh30_w141_7 :  std_logic;
signal CompressorIn_bh30_349_567 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_349_568 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_349_349 :  std_logic_vector(2 downto 0);
signal heap_bh30_w141_8 :  std_logic;
signal heap_bh30_w142_6 :  std_logic;
signal heap_bh30_w143_7 :  std_logic;
signal CompressorIn_bh30_350_569 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_350_570 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_350_350 :  std_logic_vector(2 downto 0);
signal heap_bh30_w143_8 :  std_logic;
signal heap_bh30_w144_6 :  std_logic;
signal heap_bh30_w145_7 :  std_logic;
signal CompressorIn_bh30_351_571 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_351_572 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_351_351 :  std_logic_vector(2 downto 0);
signal heap_bh30_w145_8 :  std_logic;
signal heap_bh30_w146_4 :  std_logic;
signal heap_bh30_w147_5 :  std_logic;
signal CompressorIn_bh30_352_573 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_352_574 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_352_352 :  std_logic_vector(2 downto 0);
signal heap_bh30_w157_3 :  std_logic;
signal heap_bh30_w158_2 :  std_logic;
signal heap_bh30_w159_2 :  std_logic;
signal CompressorIn_bh30_353_575 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_353_576 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_353_353 :  std_logic_vector(2 downto 0);
signal heap_bh30_w14_9 :  std_logic;
signal heap_bh30_w15_10 :  std_logic;
signal heap_bh30_w16_11 :  std_logic;
signal CompressorIn_bh30_354_577 :  std_logic_vector(2 downto 0);
signal CompressorOut_bh30_354_354 :  std_logic_vector(1 downto 0);
signal heap_bh30_w36_16 :  std_logic;
signal heap_bh30_w37_16 :  std_logic;
signal CompressorIn_bh30_355_578 :  std_logic_vector(2 downto 0);
signal CompressorOut_bh30_355_355 :  std_logic_vector(1 downto 0);
signal heap_bh30_w39_16 :  std_logic;
signal heap_bh30_w40_16 :  std_logic;
signal CompressorIn_bh30_356_579 :  std_logic_vector(2 downto 0);
signal CompressorOut_bh30_356_356 :  std_logic_vector(1 downto 0);
signal heap_bh30_w42_16 :  std_logic;
signal heap_bh30_w43_16 :  std_logic;
signal CompressorIn_bh30_357_580 :  std_logic_vector(2 downto 0);
signal CompressorOut_bh30_357_357 :  std_logic_vector(1 downto 0);
signal heap_bh30_w47_16 :  std_logic;
signal heap_bh30_w48_17 :  std_logic;
signal CompressorIn_bh30_358_581 :  std_logic_vector(2 downto 0);
signal CompressorOut_bh30_358_358 :  std_logic_vector(1 downto 0);
signal heap_bh30_w52_19 :  std_logic;
signal heap_bh30_w53_18 :  std_logic;
signal CompressorIn_bh30_359_582 :  std_logic_vector(2 downto 0);
signal CompressorOut_bh30_359_359 :  std_logic_vector(1 downto 0);
signal heap_bh30_w55_19 :  std_logic;
signal heap_bh30_w56_18 :  std_logic;
signal CompressorIn_bh30_360_583 :  std_logic_vector(2 downto 0);
signal CompressorOut_bh30_360_360 :  std_logic_vector(1 downto 0);
signal heap_bh30_w58_19 :  std_logic;
signal heap_bh30_w59_18 :  std_logic;
signal CompressorIn_bh30_361_584 :  std_logic_vector(2 downto 0);
signal CompressorOut_bh30_361_361 :  std_logic_vector(1 downto 0);
signal heap_bh30_w61_19 :  std_logic;
signal heap_bh30_w62_18 :  std_logic;
signal CompressorIn_bh30_362_585 :  std_logic_vector(2 downto 0);
signal CompressorOut_bh30_362_362 :  std_logic_vector(1 downto 0);
signal heap_bh30_w64_19 :  std_logic;
signal heap_bh30_w65_18 :  std_logic;
signal CompressorIn_bh30_363_586 :  std_logic_vector(2 downto 0);
signal CompressorOut_bh30_363_363 :  std_logic_vector(1 downto 0);
signal heap_bh30_w69_21 :  std_logic;
signal heap_bh30_w70_21 :  std_logic;
signal CompressorIn_bh30_364_587 :  std_logic_vector(2 downto 0);
signal CompressorOut_bh30_364_364 :  std_logic_vector(1 downto 0);
signal heap_bh30_w108_12 :  std_logic;
signal heap_bh30_w109_12 :  std_logic;
signal CompressorIn_bh30_365_588 :  std_logic_vector(2 downto 0);
signal CompressorOut_bh30_365_365 :  std_logic_vector(1 downto 0);
signal heap_bh30_w110_11 :  std_logic;
signal heap_bh30_w111_12 :  std_logic;
signal CompressorIn_bh30_366_589 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_366_590 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_366_366 :  std_logic_vector(2 downto 0);
signal heap_bh30_w74_23 :  std_logic;
signal heap_bh30_w75_24 :  std_logic;
signal heap_bh30_w76_23 :  std_logic;
signal CompressorIn_bh30_367_591 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_367_592 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_367_367 :  std_logic_vector(2 downto 0);
signal heap_bh30_w77_23 :  std_logic;
signal heap_bh30_w78_24 :  std_logic;
signal heap_bh30_w79_23 :  std_logic;
signal CompressorIn_bh30_368_593 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_368_594 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_368_368 :  std_logic_vector(2 downto 0);
signal heap_bh30_w80_23 :  std_logic;
signal heap_bh30_w81_24 :  std_logic;
signal heap_bh30_w82_23 :  std_logic;
signal CompressorIn_bh30_369_595 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_369_596 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_369_369 :  std_logic_vector(2 downto 0);
signal heap_bh30_w83_23 :  std_logic;
signal heap_bh30_w84_24 :  std_logic;
signal heap_bh30_w85_23 :  std_logic;
signal CompressorIn_bh30_370_597 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_370_598 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_370_370 :  std_logic_vector(2 downto 0);
signal heap_bh30_w86_23 :  std_logic;
signal heap_bh30_w87_24 :  std_logic;
signal heap_bh30_w88_23 :  std_logic;
signal CompressorIn_bh30_371_599 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_371_600 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_371_371 :  std_logic_vector(2 downto 0);
signal heap_bh30_w89_23 :  std_logic;
signal heap_bh30_w90_23 :  std_logic;
signal heap_bh30_w91_21 :  std_logic;
signal CompressorIn_bh30_372_601 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_372_602 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_372_372 :  std_logic_vector(2 downto 0);
signal heap_bh30_w92_19 :  std_logic;
signal heap_bh30_w93_18 :  std_logic;
signal heap_bh30_w94_16 :  std_logic;
signal CompressorIn_bh30_373_603 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_373_604 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_373_373 :  std_logic_vector(2 downto 0);
signal heap_bh30_w96_14 :  std_logic;
signal heap_bh30_w97_14 :  std_logic;
signal heap_bh30_w98_14 :  std_logic;
signal CompressorIn_bh30_374_605 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_374_606 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_374_374 :  std_logic_vector(2 downto 0);
signal heap_bh30_w10_10 :  std_logic;
signal heap_bh30_w11_8 :  std_logic;
signal heap_bh30_w12_10 :  std_logic;
signal CompressorIn_bh30_375_607 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_375_608 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_375_375 :  std_logic_vector(2 downto 0);
signal heap_bh30_w16_12 :  std_logic;
signal heap_bh30_w17_11 :  std_logic;
signal heap_bh30_w18_12 :  std_logic;
signal CompressorIn_bh30_376_609 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_376_610 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_376_376 :  std_logic_vector(2 downto 0);
signal heap_bh30_w35_15 :  std_logic;
signal heap_bh30_w36_17 :  std_logic;
signal heap_bh30_w37_17 :  std_logic;
signal CompressorIn_bh30_377_611 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_377_612 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_377_377 :  std_logic_vector(2 downto 0);
signal heap_bh30_w38_15 :  std_logic;
signal heap_bh30_w39_17 :  std_logic;
signal heap_bh30_w40_17 :  std_logic;
signal CompressorIn_bh30_378_613 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_378_614 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_378_378 :  std_logic_vector(2 downto 0);
signal heap_bh30_w41_15 :  std_logic;
signal heap_bh30_w42_17 :  std_logic;
signal heap_bh30_w43_17 :  std_logic;
signal CompressorIn_bh30_379_615 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_379_616 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_379_379 :  std_logic_vector(2 downto 0);
signal heap_bh30_w44_15 :  std_logic;
signal heap_bh30_w45_17 :  std_logic;
signal heap_bh30_w46_16 :  std_logic;
signal CompressorIn_bh30_380_617 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_380_618 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_380_380 :  std_logic_vector(2 downto 0);
signal heap_bh30_w49_17 :  std_logic;
signal heap_bh30_w50_18 :  std_logic;
signal heap_bh30_w51_19 :  std_logic;
signal CompressorIn_bh30_381_619 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_381_620 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_381_381 :  std_logic_vector(2 downto 0);
signal heap_bh30_w52_20 :  std_logic;
signal heap_bh30_w53_19 :  std_logic;
signal heap_bh30_w54_19 :  std_logic;
signal CompressorIn_bh30_382_621 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_382_622 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_382_382 :  std_logic_vector(2 downto 0);
signal heap_bh30_w55_20 :  std_logic;
signal heap_bh30_w56_19 :  std_logic;
signal heap_bh30_w57_19 :  std_logic;
signal CompressorIn_bh30_383_623 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_383_624 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_383_383 :  std_logic_vector(2 downto 0);
signal heap_bh30_w58_20 :  std_logic;
signal heap_bh30_w59_19 :  std_logic;
signal heap_bh30_w60_19 :  std_logic;
signal CompressorIn_bh30_384_625 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_384_626 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_384_384 :  std_logic_vector(2 downto 0);
signal heap_bh30_w61_20 :  std_logic;
signal heap_bh30_w62_19 :  std_logic;
signal heap_bh30_w63_19 :  std_logic;
signal CompressorIn_bh30_385_627 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_385_628 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_385_385 :  std_logic_vector(2 downto 0);
signal heap_bh30_w64_20 :  std_logic;
signal heap_bh30_w65_19 :  std_logic;
signal heap_bh30_w66_19 :  std_logic;
signal CompressorIn_bh30_386_629 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_386_630 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_386_386 :  std_logic_vector(2 downto 0);
signal heap_bh30_w67_21 :  std_logic;
signal heap_bh30_w68_20 :  std_logic;
signal heap_bh30_w69_22 :  std_logic;
signal CompressorIn_bh30_387_631 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_387_632 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_387_387 :  std_logic_vector(2 downto 0);
signal heap_bh30_w69_23 :  std_logic;
signal heap_bh30_w70_22 :  std_logic;
signal heap_bh30_w71_22 :  std_logic;
signal CompressorIn_bh30_388_633 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_388_634 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_388_388 :  std_logic_vector(2 downto 0);
signal heap_bh30_w72_24 :  std_logic;
signal heap_bh30_w73_23 :  std_logic;
signal heap_bh30_w74_24 :  std_logic;
signal CompressorIn_bh30_389_635 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_389_636 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_389_389 :  std_logic_vector(2 downto 0);
signal heap_bh30_w94_17 :  std_logic;
signal heap_bh30_w95_15 :  std_logic;
signal heap_bh30_w96_15 :  std_logic;
signal CompressorIn_bh30_390_637 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_390_638 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_390_390 :  std_logic_vector(2 downto 0);
signal heap_bh30_w98_15 :  std_logic;
signal heap_bh30_w99_14 :  std_logic;
signal heap_bh30_w100_14 :  std_logic;
signal CompressorIn_bh30_391_639 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_391_640 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_391_391 :  std_logic_vector(2 downto 0);
signal heap_bh30_w100_15 :  std_logic;
signal heap_bh30_w101_14 :  std_logic;
signal heap_bh30_w102_14 :  std_logic;
signal CompressorIn_bh30_392_641 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_392_642 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_392_392 :  std_logic_vector(2 downto 0);
signal heap_bh30_w102_15 :  std_logic;
signal heap_bh30_w103_14 :  std_logic;
signal heap_bh30_w104_14 :  std_logic;
signal CompressorIn_bh30_393_643 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_393_644 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_393_393 :  std_logic_vector(2 downto 0);
signal heap_bh30_w104_15 :  std_logic;
signal heap_bh30_w105_14 :  std_logic;
signal heap_bh30_w106_14 :  std_logic;
signal CompressorIn_bh30_394_645 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_394_646 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_394_394 :  std_logic_vector(2 downto 0);
signal heap_bh30_w106_15 :  std_logic;
signal heap_bh30_w107_14 :  std_logic;
signal heap_bh30_w108_13 :  std_logic;
signal CompressorIn_bh30_395_647 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_395_648 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_395_395 :  std_logic_vector(2 downto 0);
signal heap_bh30_w108_14 :  std_logic;
signal heap_bh30_w109_13 :  std_logic;
signal heap_bh30_w110_12 :  std_logic;
signal CompressorIn_bh30_396_649 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_396_650 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_396_396 :  std_logic_vector(2 downto 0);
signal heap_bh30_w111_13 :  std_logic;
signal heap_bh30_w112_10 :  std_logic;
signal heap_bh30_w113_11 :  std_logic;
signal CompressorIn_bh30_397_651 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_397_652 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_397_397 :  std_logic_vector(2 downto 0);
signal heap_bh30_w130_9 :  std_logic;
signal heap_bh30_w131_10 :  std_logic;
signal heap_bh30_w132_8 :  std_logic;
signal CompressorIn_bh30_398_653 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_398_654 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_398_398 :  std_logic_vector(2 downto 0);
signal heap_bh30_w147_6 :  std_logic;
signal heap_bh30_w148_4 :  std_logic;
signal heap_bh30_w149_5 :  std_logic;
signal CompressorIn_bh30_399_655 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_399_656 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_399_399 :  std_logic_vector(2 downto 0);
signal heap_bh30_w159_3 :  std_logic;
signal heap_bh30_w160_2 :  std_logic;
signal heap_bh30_w161_2 :  std_logic;
signal CompressorIn_bh30_400_657 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_400_658 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_400_400 :  std_logic_vector(2 downto 0);
signal heap_bh30_w21_13 :  std_logic;
signal heap_bh30_w22_12 :  std_logic;
signal heap_bh30_w23_13 :  std_logic;
signal CompressorIn_bh30_401_659 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_401_660 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_401_401 :  std_logic_vector(2 downto 0);
signal heap_bh30_w24_14 :  std_logic;
signal heap_bh30_w25_15 :  std_logic;
signal heap_bh30_w26_14 :  std_logic;
signal CompressorIn_bh30_402_661 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_402_662 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_402_402 :  std_logic_vector(2 downto 0);
signal heap_bh30_w27_14 :  std_logic;
signal heap_bh30_w28_15 :  std_logic;
signal heap_bh30_w29_14 :  std_logic;
signal CompressorIn_bh30_403_663 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_403_664 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_403_403 :  std_logic_vector(2 downto 0);
signal heap_bh30_w30_14 :  std_logic;
signal heap_bh30_w31_15 :  std_logic;
signal heap_bh30_w32_14 :  std_logic;
signal CompressorIn_bh30_404_665 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_404_666 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_404_404 :  std_logic_vector(2 downto 0);
signal heap_bh30_w33_15 :  std_logic;
signal heap_bh30_w34_16 :  std_logic;
signal heap_bh30_w35_16 :  std_logic;
signal CompressorIn_bh30_405_667 :  std_logic_vector(2 downto 0);
signal CompressorOut_bh30_405_405 :  std_logic_vector(1 downto 0);
signal heap_bh30_w76_24 :  std_logic;
signal heap_bh30_w77_24 :  std_logic;
signal CompressorIn_bh30_406_668 :  std_logic_vector(2 downto 0);
signal CompressorOut_bh30_406_406 :  std_logic_vector(1 downto 0);
signal heap_bh30_w79_24 :  std_logic;
signal heap_bh30_w80_24 :  std_logic;
signal CompressorIn_bh30_407_669 :  std_logic_vector(2 downto 0);
signal CompressorOut_bh30_407_407 :  std_logic_vector(1 downto 0);
signal heap_bh30_w82_24 :  std_logic;
signal heap_bh30_w83_24 :  std_logic;
signal CompressorIn_bh30_408_670 :  std_logic_vector(2 downto 0);
signal CompressorOut_bh30_408_408 :  std_logic_vector(1 downto 0);
signal heap_bh30_w85_24 :  std_logic;
signal heap_bh30_w86_24 :  std_logic;
signal CompressorIn_bh30_409_671 :  std_logic_vector(2 downto 0);
signal CompressorOut_bh30_409_409 :  std_logic_vector(1 downto 0);
signal heap_bh30_w88_24 :  std_logic;
signal heap_bh30_w89_24 :  std_logic;
signal CompressorIn_bh30_410_672 :  std_logic_vector(2 downto 0);
signal CompressorOut_bh30_410_410 :  std_logic_vector(1 downto 0);
signal heap_bh30_w91_22 :  std_logic;
signal heap_bh30_w92_20 :  std_logic;
signal CompressorIn_bh30_411_673 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_411_674 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_411_411 :  std_logic_vector(2 downto 0);
signal heap_bh30_w46_17 :  std_logic;
signal heap_bh30_w47_17 :  std_logic;
signal heap_bh30_w48_18 :  std_logic;
signal CompressorIn_bh30_412_675 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_412_676 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_412_412 :  std_logic_vector(2 downto 0);
signal heap_bh30_w75_25 :  std_logic;
signal heap_bh30_w76_25 :  std_logic;
signal heap_bh30_w77_25 :  std_logic;
signal CompressorIn_bh30_413_677 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_413_678 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_413_413 :  std_logic_vector(2 downto 0);
signal heap_bh30_w78_25 :  std_logic;
signal heap_bh30_w79_25 :  std_logic;
signal heap_bh30_w80_25 :  std_logic;
signal CompressorIn_bh30_414_679 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_414_680 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_414_414 :  std_logic_vector(2 downto 0);
signal heap_bh30_w81_25 :  std_logic;
signal heap_bh30_w82_25 :  std_logic;
signal heap_bh30_w83_25 :  std_logic;
signal CompressorIn_bh30_415_681 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_415_682 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_415_415 :  std_logic_vector(2 downto 0);
signal heap_bh30_w84_25 :  std_logic;
signal heap_bh30_w85_25 :  std_logic;
signal heap_bh30_w86_25 :  std_logic;
signal CompressorIn_bh30_416_683 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_416_684 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_416_416 :  std_logic_vector(2 downto 0);
signal heap_bh30_w87_25 :  std_logic;
signal heap_bh30_w88_25 :  std_logic;
signal heap_bh30_w89_25 :  std_logic;
signal CompressorIn_bh30_417_685 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_417_686 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_417_417 :  std_logic_vector(2 downto 0);
signal heap_bh30_w90_24 :  std_logic;
signal heap_bh30_w91_23 :  std_logic;
signal heap_bh30_w92_21 :  std_logic;
signal CompressorIn_bh30_418_687 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_418_688 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_418_418 :  std_logic_vector(2 downto 0);
signal heap_bh30_w93_19 :  std_logic;
signal heap_bh30_w94_18 :  std_logic;
signal heap_bh30_w95_16 :  std_logic;
signal CompressorIn_bh30_419_689 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_419_690 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_419_419 :  std_logic_vector(2 downto 0);
signal heap_bh30_w97_15 :  std_logic;
signal heap_bh30_w98_16 :  std_logic;
signal heap_bh30_w99_15 :  std_logic;
signal CompressorIn_bh30_420_691 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_420_692 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_420_420 :  std_logic_vector(2 downto 0);
signal heap_bh30_w113_12 :  std_logic;
signal heap_bh30_w114_10 :  std_logic;
signal heap_bh30_w115_11 :  std_logic;
signal CompressorIn_bh30_421_693 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_421_694 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_421_421 :  std_logic_vector(2 downto 0);
signal heap_bh30_w132_9 :  std_logic;
signal heap_bh30_w133_9 :  std_logic;
signal heap_bh30_w134_7 :  std_logic;
signal CompressorIn_bh30_422_695 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_422_696 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_422_422 :  std_logic_vector(2 downto 0);
signal heap_bh30_w149_6 :  std_logic;
signal heap_bh30_w150_4 :  std_logic;
signal heap_bh30_w151_5 :  std_logic;
signal CompressorIn_bh30_423_697 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_423_698 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_423_423 :  std_logic_vector(2 downto 0);
signal heap_bh30_w161_3 :  std_logic;
signal heap_bh30_w162_2 :  std_logic;
signal heap_bh30_w163_1 :  std_logic;
signal CompressorIn_bh30_424_699 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_424_700 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_424_424 :  std_logic_vector(2 downto 0);
signal heap_bh30_w18_13 :  std_logic;
signal heap_bh30_w19_12 :  std_logic;
signal heap_bh30_w20_12 :  std_logic;
signal CompressorIn_bh30_425_701 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_425_702 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_425_425 :  std_logic_vector(2 downto 0);
signal heap_bh30_w26_15 :  std_logic;
signal heap_bh30_w27_15 :  std_logic;
signal heap_bh30_w28_16 :  std_logic;
signal CompressorIn_bh30_426_703 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_426_704 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_426_426 :  std_logic_vector(2 downto 0);
signal heap_bh30_w29_15 :  std_logic;
signal heap_bh30_w30_15 :  std_logic;
signal heap_bh30_w31_16 :  std_logic;
signal CompressorIn_bh30_427_705 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_427_706 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_427_427 :  std_logic_vector(2 downto 0);
signal heap_bh30_w32_15 :  std_logic;
signal heap_bh30_w33_16 :  std_logic;
signal heap_bh30_w34_17 :  std_logic;
signal CompressorIn_bh30_428_707 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_428_708 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_428_428 :  std_logic_vector(2 downto 0);
signal heap_bh30_w37_18 :  std_logic;
signal heap_bh30_w38_16 :  std_logic;
signal heap_bh30_w39_18 :  std_logic;
signal CompressorIn_bh30_429_709 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_429_710 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_429_429 :  std_logic_vector(2 downto 0);
signal heap_bh30_w40_18 :  std_logic;
signal heap_bh30_w41_16 :  std_logic;
signal heap_bh30_w42_18 :  std_logic;
signal CompressorIn_bh30_430_711 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_430_712 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_430_430 :  std_logic_vector(2 downto 0);
signal heap_bh30_w43_18 :  std_logic;
signal heap_bh30_w44_16 :  std_logic;
signal heap_bh30_w45_18 :  std_logic;
signal CompressorIn_bh30_431_713 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_431_714 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_431_431 :  std_logic_vector(2 downto 0);
signal heap_bh30_w51_20 :  std_logic;
signal heap_bh30_w52_21 :  std_logic;
signal heap_bh30_w53_20 :  std_logic;
signal CompressorIn_bh30_432_715 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_432_716 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_432_432 :  std_logic_vector(2 downto 0);
signal heap_bh30_w54_20 :  std_logic;
signal heap_bh30_w55_21 :  std_logic;
signal heap_bh30_w56_20 :  std_logic;
signal CompressorIn_bh30_433_717 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_433_718 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_433_433 :  std_logic_vector(2 downto 0);
signal heap_bh30_w57_20 :  std_logic;
signal heap_bh30_w58_21 :  std_logic;
signal heap_bh30_w59_20 :  std_logic;
signal CompressorIn_bh30_434_719 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_434_720 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_434_434 :  std_logic_vector(2 downto 0);
signal heap_bh30_w60_20 :  std_logic;
signal heap_bh30_w61_21 :  std_logic;
signal heap_bh30_w62_20 :  std_logic;
signal CompressorIn_bh30_435_721 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_435_722 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_435_435 :  std_logic_vector(2 downto 0);
signal heap_bh30_w63_20 :  std_logic;
signal heap_bh30_w64_21 :  std_logic;
signal heap_bh30_w65_20 :  std_logic;
signal CompressorIn_bh30_436_723 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_436_724 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_436_436 :  std_logic_vector(2 downto 0);
signal heap_bh30_w66_20 :  std_logic;
signal heap_bh30_w67_22 :  std_logic;
signal heap_bh30_w68_21 :  std_logic;
signal CompressorIn_bh30_437_725 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_437_726 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_437_437 :  std_logic_vector(2 downto 0);
signal heap_bh30_w71_23 :  std_logic;
signal heap_bh30_w72_25 :  std_logic;
signal heap_bh30_w73_24 :  std_logic;
signal CompressorIn_bh30_438_727 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_438_728 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_438_438 :  std_logic_vector(2 downto 0);
signal heap_bh30_w110_13 :  std_logic;
signal heap_bh30_w111_14 :  std_logic;
signal heap_bh30_w112_11 :  std_logic;
signal CompressorIn_bh30_439_729 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_439_730 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_439_439 :  std_logic_vector(2 downto 0);
signal heap_bh30_w68_22 :  std_logic;
signal heap_bh30_w69_24 :  std_logic;
signal heap_bh30_w70_23 :  std_logic;
signal CompressorIn_bh30_440_731 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_440_732 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_440_440 :  std_logic_vector(2 downto 0);
signal heap_bh30_w73_25 :  std_logic;
signal heap_bh30_w74_25 :  std_logic;
signal heap_bh30_w75_26 :  std_logic;
signal CompressorIn_bh30_441_733 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_441_734 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_441_441 :  std_logic_vector(2 downto 0);
signal heap_bh30_w95_17 :  std_logic;
signal heap_bh30_w96_16 :  std_logic;
signal heap_bh30_w97_16 :  std_logic;
signal CompressorIn_bh30_442_735 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_442_736 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_442_442 :  std_logic_vector(2 downto 0);
signal heap_bh30_w99_16 :  std_logic;
signal heap_bh30_w100_16 :  std_logic;
signal heap_bh30_w101_15 :  std_logic;
signal CompressorIn_bh30_443_737 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_443_738 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_443_443 :  std_logic_vector(2 downto 0);
signal heap_bh30_w115_12 :  std_logic;
signal heap_bh30_w116_10 :  std_logic;
signal heap_bh30_w117_11 :  std_logic;
signal CompressorIn_bh30_444_739 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_444_740 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_444_444 :  std_logic_vector(2 downto 0);
signal heap_bh30_w151_6 :  std_logic;
signal heap_bh30_w152_4 :  std_logic;
signal heap_bh30_w153_5 :  std_logic;
signal CompressorIn_bh30_445_741 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_445_742 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_445_445 :  std_logic_vector(2 downto 0);
signal heap_bh30_w48_19 :  std_logic;
signal heap_bh30_w49_18 :  std_logic;
signal heap_bh30_w50_19 :  std_logic;
signal CompressorIn_bh30_446_743 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_446_744 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_446_446 :  std_logic_vector(2 downto 0);
signal heap_bh30_w53_21 :  std_logic;
signal heap_bh30_w54_21 :  std_logic;
signal heap_bh30_w55_22 :  std_logic;
signal CompressorIn_bh30_447_745 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_447_746 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_447_447 :  std_logic_vector(2 downto 0);
signal heap_bh30_w56_21 :  std_logic;
signal heap_bh30_w57_21 :  std_logic;
signal heap_bh30_w58_22 :  std_logic;
signal CompressorIn_bh30_448_747 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_448_748 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_448_448 :  std_logic_vector(2 downto 0);
signal heap_bh30_w59_21 :  std_logic;
signal heap_bh30_w60_21 :  std_logic;
signal heap_bh30_w61_22 :  std_logic;
signal CompressorIn_bh30_449_749 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_449_750 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_449_449 :  std_logic_vector(2 downto 0);
signal heap_bh30_w62_21 :  std_logic;
signal heap_bh30_w63_21 :  std_logic;
signal heap_bh30_w64_22 :  std_logic;
signal CompressorIn_bh30_450_751 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_450_752 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_450_450 :  std_logic_vector(2 downto 0);
signal heap_bh30_w65_21 :  std_logic;
signal heap_bh30_w66_21 :  std_logic;
signal heap_bh30_w67_23 :  std_logic;
signal CompressorIn_bh30_451_753 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_451_754 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_451_451 :  std_logic_vector(2 downto 0);
signal heap_bh30_w77_26 :  std_logic;
signal heap_bh30_w78_26 :  std_logic;
signal heap_bh30_w79_26 :  std_logic;
signal CompressorIn_bh30_452_755 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_452_756 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_452_452 :  std_logic_vector(2 downto 0);
signal heap_bh30_w80_26 :  std_logic;
signal heap_bh30_w81_26 :  std_logic;
signal heap_bh30_w82_26 :  std_logic;
signal CompressorIn_bh30_453_757 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_453_758 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_453_453 :  std_logic_vector(2 downto 0);
signal heap_bh30_w83_26 :  std_logic;
signal heap_bh30_w84_26 :  std_logic;
signal heap_bh30_w85_26 :  std_logic;
signal CompressorIn_bh30_454_759 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_454_760 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_454_454 :  std_logic_vector(2 downto 0);
signal heap_bh30_w86_26 :  std_logic;
signal heap_bh30_w87_26 :  std_logic;
signal heap_bh30_w88_26 :  std_logic;
signal CompressorIn_bh30_455_761 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_455_762 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_455_455 :  std_logic_vector(2 downto 0);
signal heap_bh30_w89_26 :  std_logic;
signal heap_bh30_w90_25 :  std_logic;
signal heap_bh30_w91_24 :  std_logic;
signal CompressorIn_bh30_456_763 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_456_764 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_456_456 :  std_logic_vector(2 downto 0);
signal heap_bh30_w92_22 :  std_logic;
signal heap_bh30_w93_20 :  std_logic;
signal heap_bh30_w94_19 :  std_logic;
signal CompressorIn_bh30_457_765 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_457_766 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_457_457 :  std_logic_vector(2 downto 0);
signal heap_bh30_w112_12 :  std_logic;
signal heap_bh30_w113_13 :  std_logic;
signal heap_bh30_w114_11 :  std_logic;
signal CompressorIn_bh30_458_767 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_458_768 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_458_458 :  std_logic_vector(2 downto 0);
signal heap_bh30_w101_16 :  std_logic;
signal heap_bh30_w102_16 :  std_logic;
signal heap_bh30_w103_15 :  std_logic;
signal CompressorIn_bh30_459_769 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_459_770 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_459_459 :  std_logic_vector(2 downto 0);
signal heap_bh30_w117_12 :  std_logic;
signal heap_bh30_w118_10 :  std_logic;
signal heap_bh30_w119_11 :  std_logic;
signal CompressorIn_bh30_460_771 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_460_772 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_460_460 :  std_logic_vector(2 downto 0);
signal heap_bh30_w153_6 :  std_logic;
signal heap_bh30_w154_4 :  std_logic;
signal heap_bh30_w155_5 :  std_logic;
signal CompressorIn_bh30_461_773 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_461_774 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_461_461 :  std_logic_vector(2 downto 0);
signal heap_bh30_w70_24 :  std_logic;
signal heap_bh30_w71_24 :  std_logic;
signal heap_bh30_w72_26 :  std_logic;
signal CompressorIn_bh30_462_775 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_462_776 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_462_462 :  std_logic_vector(2 downto 0);
signal heap_bh30_w103_16 :  std_logic;
signal heap_bh30_w104_16 :  std_logic;
signal heap_bh30_w105_15 :  std_logic;
signal CompressorIn_bh30_463_777 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_463_778 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_463_463 :  std_logic_vector(2 downto 0);
signal heap_bh30_w119_12 :  std_logic;
signal heap_bh30_w120_10 :  std_logic;
signal heap_bh30_w121_11 :  std_logic;
signal CompressorIn_bh30_464_779 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_464_780 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_464_464 :  std_logic_vector(2 downto 0);
signal heap_bh30_w155_6 :  std_logic;
signal heap_bh30_w156_3 :  std_logic;
signal heap_bh30_w157_4 :  std_logic;
signal CompressorIn_bh30_465_781 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_465_782 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_465_465 :  std_logic_vector(2 downto 0);
signal heap_bh30_w105_16 :  std_logic;
signal heap_bh30_w106_16 :  std_logic;
signal heap_bh30_w107_15 :  std_logic;
signal CompressorIn_bh30_466_783 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_466_784 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_466_466 :  std_logic_vector(2 downto 0);
signal heap_bh30_w121_12 :  std_logic;
signal heap_bh30_w122_10 :  std_logic;
signal heap_bh30_w123_11 :  std_logic;
signal CompressorIn_bh30_467_785 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_467_786 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_467_467 :  std_logic_vector(2 downto 0);
signal heap_bh30_w107_16 :  std_logic;
signal heap_bh30_w108_15 :  std_logic;
signal heap_bh30_w109_14 :  std_logic;
signal CompressorIn_bh30_468_787 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_468_788 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_468_468 :  std_logic_vector(2 downto 0);
signal heap_bh30_w123_12 :  std_logic;
signal heap_bh30_w124_10 :  std_logic;
signal heap_bh30_w125_11 :  std_logic;
signal CompressorIn_bh30_469_789 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_469_790 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_469_469 :  std_logic_vector(2 downto 0);
signal heap_bh30_w125_12 :  std_logic;
signal heap_bh30_w126_10 :  std_logic;
signal heap_bh30_w127_11 :  std_logic;
signal CompressorIn_bh30_470_791 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_470_792 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_470_470 :  std_logic_vector(2 downto 0);
signal heap_bh30_w109_15 :  std_logic;
signal heap_bh30_w110_14 :  std_logic;
signal heap_bh30_w111_15 :  std_logic;
signal CompressorIn_bh30_471_793 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_471_794 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_471_471 :  std_logic_vector(2 downto 0);
signal heap_bh30_w127_12 :  std_logic;
signal heap_bh30_w128_10 :  std_logic;
signal heap_bh30_w129_10 :  std_logic;
signal CompressorIn_bh30_472_795 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_472_796 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_472_472 :  std_logic_vector(2 downto 0);
signal heap_bh30_w129_11 :  std_logic;
signal heap_bh30_w130_10 :  std_logic;
signal heap_bh30_w131_11 :  std_logic;
signal finalAdderIn0_bh30 :  std_logic_vector(180 downto 0);
signal finalAdderIn1_bh30 :  std_logic_vector(180 downto 0);
signal finalAdderCin_bh30 :  std_logic;
signal finalAdderOut_bh30 :  std_logic_vector(180 downto 0);
signal CompressionResult30 :  std_logic_vector(180 downto 0);
attribute rom_extract: string;
attribute rom_style: string;
attribute rom_extract of SmallMultTableP3x3r6XuYu_comb_uid103: component is "yes";
attribute rom_extract of SmallMultTableP3x3r6XuYu_comb_uid138: component is "yes";
attribute rom_extract of SmallMultTableP3x3r6XuYu_comb_uid33: component is "yes";
attribute rom_extract of SmallMultTableP3x3r6XuYu_comb_uid68: component is "yes";
attribute rom_style of SmallMultTableP3x3r6XuYu_comb_uid103: component is "distributed";
attribute rom_style of SmallMultTableP3x3r6XuYu_comb_uid138: component is "distributed";
attribute rom_style of SmallMultTableP3x3r6XuYu_comb_uid33: component is "distributed";
attribute rom_style of SmallMultTableP3x3r6XuYu_comb_uid68: component is "distributed";
begin
   XX_m29 <= X ;
   YY_m29 <= Y ;
   -- code generated by IntMultiplier::buildHeapLogicOnly()
   -- buildheaplogiconly called for lsbX=66 lsbY=0 msbX=90 msbY=5
   Xp_m29b31 <= XX_m29(89 downto 66) & "";
   Yp_m29b31 <= YY_m29(4 downto 0) & "0";
   x_m29b31_0 <= Xp_m29b31(2 downto 0);
   x_m29b31_1 <= Xp_m29b31(5 downto 3);
   x_m29b31_2 <= Xp_m29b31(8 downto 6);
   x_m29b31_3 <= Xp_m29b31(11 downto 9);
   x_m29b31_4 <= Xp_m29b31(14 downto 12);
   x_m29b31_5 <= Xp_m29b31(17 downto 15);
   x_m29b31_6 <= Xp_m29b31(20 downto 18);
   x_m29b31_7 <= Xp_m29b31(23 downto 21);
   y_m29b31_0 <= Yp_m29b31(2 downto 0);
   y_m29b31_1 <= Yp_m29b31(5 downto 3);
   -- Partial product row number 0
   Y0X0_31_m29 <= y_m29b31_0 & x_m29b31_0;
   PP_m29_31X0Y0_Tbl: SmallMultTableP3x3r6XuYu_comb_uid33
      port map ( X => Y0X0_31_m29,
                 Y => PP31X0Y0_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w66_0 <= PP31X0Y0_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w67_0 <= PP31X0Y0_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w68_0 <= PP31X0Y0_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w69_0 <= PP31X0Y0_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w70_0 <= PP31X0Y0_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y0X1_31_m29 <= y_m29b31_0 & x_m29b31_1;
   PP_m29_31X1Y0_Tbl: SmallMultTableP3x3r6XuYu_comb_uid33
      port map ( X => Y0X1_31_m29,
                 Y => PP31X1Y0_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w69_1 <= PP31X1Y0_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w70_1 <= PP31X1Y0_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w71_0 <= PP31X1Y0_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w72_0 <= PP31X1Y0_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w73_0 <= PP31X1Y0_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y0X2_31_m29 <= y_m29b31_0 & x_m29b31_2;
   PP_m29_31X2Y0_Tbl: SmallMultTableP3x3r6XuYu_comb_uid33
      port map ( X => Y0X2_31_m29,
                 Y => PP31X2Y0_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w72_1 <= PP31X2Y0_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w73_1 <= PP31X2Y0_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w74_0 <= PP31X2Y0_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w75_0 <= PP31X2Y0_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w76_0 <= PP31X2Y0_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y0X3_31_m29 <= y_m29b31_0 & x_m29b31_3;
   PP_m29_31X3Y0_Tbl: SmallMultTableP3x3r6XuYu_comb_uid33
      port map ( X => Y0X3_31_m29,
                 Y => PP31X3Y0_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w75_1 <= PP31X3Y0_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w76_1 <= PP31X3Y0_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w77_0 <= PP31X3Y0_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w78_0 <= PP31X3Y0_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w79_0 <= PP31X3Y0_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y0X4_31_m29 <= y_m29b31_0 & x_m29b31_4;
   PP_m29_31X4Y0_Tbl: SmallMultTableP3x3r6XuYu_comb_uid33
      port map ( X => Y0X4_31_m29,
                 Y => PP31X4Y0_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w78_1 <= PP31X4Y0_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w79_1 <= PP31X4Y0_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w80_0 <= PP31X4Y0_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w81_0 <= PP31X4Y0_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w82_0 <= PP31X4Y0_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y0X5_31_m29 <= y_m29b31_0 & x_m29b31_5;
   PP_m29_31X5Y0_Tbl: SmallMultTableP3x3r6XuYu_comb_uid33
      port map ( X => Y0X5_31_m29,
                 Y => PP31X5Y0_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w81_1 <= PP31X5Y0_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w82_1 <= PP31X5Y0_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w83_0 <= PP31X5Y0_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w84_0 <= PP31X5Y0_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w85_0 <= PP31X5Y0_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y0X6_31_m29 <= y_m29b31_0 & x_m29b31_6;
   PP_m29_31X6Y0_Tbl: SmallMultTableP3x3r6XuYu_comb_uid33
      port map ( X => Y0X6_31_m29,
                 Y => PP31X6Y0_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w84_1 <= PP31X6Y0_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w85_1 <= PP31X6Y0_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w86_0 <= PP31X6Y0_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w87_0 <= PP31X6Y0_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w88_0 <= PP31X6Y0_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y0X7_31_m29 <= y_m29b31_0 & x_m29b31_7;
   PP_m29_31X7Y0_Tbl: SmallMultTableP3x3r6XuYu_comb_uid33
      port map ( X => Y0X7_31_m29,
                 Y => PP31X7Y0_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w87_1 <= PP31X7Y0_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w88_1 <= PP31X7Y0_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w89_0 <= PP31X7Y0_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w90_0 <= PP31X7Y0_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w91_0 <= PP31X7Y0_m29(5); -- cycle= 0 cp= 5.9176e-10

   -- Partial product row number 1
   Y1X0_31_m29 <= y_m29b31_1 & x_m29b31_0;
   PP_m29_31X0Y1_Tbl: SmallMultTableP3x3r6XuYu_comb_uid33
      port map ( X => Y1X0_31_m29,
                 Y => PP31X0Y1_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w68_1 <= PP31X0Y1_m29(0); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w69_2 <= PP31X0Y1_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w70_2 <= PP31X0Y1_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w71_1 <= PP31X0Y1_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w72_2 <= PP31X0Y1_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w73_2 <= PP31X0Y1_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y1X1_31_m29 <= y_m29b31_1 & x_m29b31_1;
   PP_m29_31X1Y1_Tbl: SmallMultTableP3x3r6XuYu_comb_uid33
      port map ( X => Y1X1_31_m29,
                 Y => PP31X1Y1_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w71_2 <= PP31X1Y1_m29(0); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w72_3 <= PP31X1Y1_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w73_3 <= PP31X1Y1_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w74_1 <= PP31X1Y1_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w75_2 <= PP31X1Y1_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w76_2 <= PP31X1Y1_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y1X2_31_m29 <= y_m29b31_1 & x_m29b31_2;
   PP_m29_31X2Y1_Tbl: SmallMultTableP3x3r6XuYu_comb_uid33
      port map ( X => Y1X2_31_m29,
                 Y => PP31X2Y1_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w74_2 <= PP31X2Y1_m29(0); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w75_3 <= PP31X2Y1_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w76_3 <= PP31X2Y1_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w77_1 <= PP31X2Y1_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w78_2 <= PP31X2Y1_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w79_2 <= PP31X2Y1_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y1X3_31_m29 <= y_m29b31_1 & x_m29b31_3;
   PP_m29_31X3Y1_Tbl: SmallMultTableP3x3r6XuYu_comb_uid33
      port map ( X => Y1X3_31_m29,
                 Y => PP31X3Y1_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w77_2 <= PP31X3Y1_m29(0); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w78_3 <= PP31X3Y1_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w79_3 <= PP31X3Y1_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w80_1 <= PP31X3Y1_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w81_2 <= PP31X3Y1_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w82_2 <= PP31X3Y1_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y1X4_31_m29 <= y_m29b31_1 & x_m29b31_4;
   PP_m29_31X4Y1_Tbl: SmallMultTableP3x3r6XuYu_comb_uid33
      port map ( X => Y1X4_31_m29,
                 Y => PP31X4Y1_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w80_2 <= PP31X4Y1_m29(0); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w81_3 <= PP31X4Y1_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w82_3 <= PP31X4Y1_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w83_1 <= PP31X4Y1_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w84_2 <= PP31X4Y1_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w85_2 <= PP31X4Y1_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y1X5_31_m29 <= y_m29b31_1 & x_m29b31_5;
   PP_m29_31X5Y1_Tbl: SmallMultTableP3x3r6XuYu_comb_uid33
      port map ( X => Y1X5_31_m29,
                 Y => PP31X5Y1_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w83_2 <= PP31X5Y1_m29(0); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w84_3 <= PP31X5Y1_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w85_3 <= PP31X5Y1_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w86_1 <= PP31X5Y1_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w87_2 <= PP31X5Y1_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w88_2 <= PP31X5Y1_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y1X6_31_m29 <= y_m29b31_1 & x_m29b31_6;
   PP_m29_31X6Y1_Tbl: SmallMultTableP3x3r6XuYu_comb_uid33
      port map ( X => Y1X6_31_m29,
                 Y => PP31X6Y1_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w86_2 <= PP31X6Y1_m29(0); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w87_3 <= PP31X6Y1_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w88_3 <= PP31X6Y1_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w89_1 <= PP31X6Y1_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w90_1 <= PP31X6Y1_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w91_1 <= PP31X6Y1_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y1X7_31_m29 <= y_m29b31_1 & x_m29b31_7;
   PP_m29_31X7Y1_Tbl: SmallMultTableP3x3r6XuYu_comb_uid33
      port map ( X => Y1X7_31_m29,
                 Y => PP31X7Y1_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w89_2 <= PP31X7Y1_m29(0); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w90_2 <= PP31X7Y1_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w91_2 <= PP31X7Y1_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w92_0 <= PP31X7Y1_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w93_0 <= PP31X7Y1_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w94_0 <= PP31X7Y1_m29(5); -- cycle= 0 cp= 5.9176e-10

   -- code generated by IntMultiplier::buildHeapLogicOnly()
   -- buildheaplogiconly called for lsbX=42 lsbY=0 msbX=66 msbY=5
   Xp_m29b66 <= XX_m29(65 downto 42) & "";
   Yp_m29b66 <= YY_m29(4 downto 0) & "0";
   x_m29b66_0 <= Xp_m29b66(2 downto 0);
   x_m29b66_1 <= Xp_m29b66(5 downto 3);
   x_m29b66_2 <= Xp_m29b66(8 downto 6);
   x_m29b66_3 <= Xp_m29b66(11 downto 9);
   x_m29b66_4 <= Xp_m29b66(14 downto 12);
   x_m29b66_5 <= Xp_m29b66(17 downto 15);
   x_m29b66_6 <= Xp_m29b66(20 downto 18);
   x_m29b66_7 <= Xp_m29b66(23 downto 21);
   y_m29b66_0 <= Yp_m29b66(2 downto 0);
   y_m29b66_1 <= Yp_m29b66(5 downto 3);
   -- Partial product row number 0
   Y0X0_66_m29 <= y_m29b66_0 & x_m29b66_0;
   PP_m29_66X0Y0_Tbl: SmallMultTableP3x3r6XuYu_comb_uid68
      port map ( X => Y0X0_66_m29,
                 Y => PP66X0Y0_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w42_0 <= PP66X0Y0_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w43_0 <= PP66X0Y0_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w44_0 <= PP66X0Y0_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w45_0 <= PP66X0Y0_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w46_0 <= PP66X0Y0_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y0X1_66_m29 <= y_m29b66_0 & x_m29b66_1;
   PP_m29_66X1Y0_Tbl: SmallMultTableP3x3r6XuYu_comb_uid68
      port map ( X => Y0X1_66_m29,
                 Y => PP66X1Y0_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w45_1 <= PP66X1Y0_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w46_1 <= PP66X1Y0_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w47_0 <= PP66X1Y0_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w48_0 <= PP66X1Y0_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w49_0 <= PP66X1Y0_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y0X2_66_m29 <= y_m29b66_0 & x_m29b66_2;
   PP_m29_66X2Y0_Tbl: SmallMultTableP3x3r6XuYu_comb_uid68
      port map ( X => Y0X2_66_m29,
                 Y => PP66X2Y0_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w48_1 <= PP66X2Y0_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w49_1 <= PP66X2Y0_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w50_0 <= PP66X2Y0_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w51_0 <= PP66X2Y0_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w52_0 <= PP66X2Y0_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y0X3_66_m29 <= y_m29b66_0 & x_m29b66_3;
   PP_m29_66X3Y0_Tbl: SmallMultTableP3x3r6XuYu_comb_uid68
      port map ( X => Y0X3_66_m29,
                 Y => PP66X3Y0_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w51_1 <= PP66X3Y0_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w52_1 <= PP66X3Y0_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w53_0 <= PP66X3Y0_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w54_0 <= PP66X3Y0_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w55_0 <= PP66X3Y0_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y0X4_66_m29 <= y_m29b66_0 & x_m29b66_4;
   PP_m29_66X4Y0_Tbl: SmallMultTableP3x3r6XuYu_comb_uid68
      port map ( X => Y0X4_66_m29,
                 Y => PP66X4Y0_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w54_1 <= PP66X4Y0_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w55_1 <= PP66X4Y0_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w56_0 <= PP66X4Y0_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w57_0 <= PP66X4Y0_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w58_0 <= PP66X4Y0_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y0X5_66_m29 <= y_m29b66_0 & x_m29b66_5;
   PP_m29_66X5Y0_Tbl: SmallMultTableP3x3r6XuYu_comb_uid68
      port map ( X => Y0X5_66_m29,
                 Y => PP66X5Y0_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w57_1 <= PP66X5Y0_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w58_1 <= PP66X5Y0_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w59_0 <= PP66X5Y0_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w60_0 <= PP66X5Y0_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w61_0 <= PP66X5Y0_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y0X6_66_m29 <= y_m29b66_0 & x_m29b66_6;
   PP_m29_66X6Y0_Tbl: SmallMultTableP3x3r6XuYu_comb_uid68
      port map ( X => Y0X6_66_m29,
                 Y => PP66X6Y0_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w60_1 <= PP66X6Y0_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w61_1 <= PP66X6Y0_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w62_0 <= PP66X6Y0_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w63_0 <= PP66X6Y0_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w64_0 <= PP66X6Y0_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y0X7_66_m29 <= y_m29b66_0 & x_m29b66_7;
   PP_m29_66X7Y0_Tbl: SmallMultTableP3x3r6XuYu_comb_uid68
      port map ( X => Y0X7_66_m29,
                 Y => PP66X7Y0_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w63_1 <= PP66X7Y0_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w64_1 <= PP66X7Y0_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w65_0 <= PP66X7Y0_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w66_1 <= PP66X7Y0_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w67_1 <= PP66X7Y0_m29(5); -- cycle= 0 cp= 5.9176e-10

   -- Partial product row number 1
   Y1X0_66_m29 <= y_m29b66_1 & x_m29b66_0;
   PP_m29_66X0Y1_Tbl: SmallMultTableP3x3r6XuYu_comb_uid68
      port map ( X => Y1X0_66_m29,
                 Y => PP66X0Y1_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w44_1 <= PP66X0Y1_m29(0); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w45_2 <= PP66X0Y1_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w46_2 <= PP66X0Y1_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w47_1 <= PP66X0Y1_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w48_2 <= PP66X0Y1_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w49_2 <= PP66X0Y1_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y1X1_66_m29 <= y_m29b66_1 & x_m29b66_1;
   PP_m29_66X1Y1_Tbl: SmallMultTableP3x3r6XuYu_comb_uid68
      port map ( X => Y1X1_66_m29,
                 Y => PP66X1Y1_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w47_2 <= PP66X1Y1_m29(0); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w48_3 <= PP66X1Y1_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w49_3 <= PP66X1Y1_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w50_1 <= PP66X1Y1_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w51_2 <= PP66X1Y1_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w52_2 <= PP66X1Y1_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y1X2_66_m29 <= y_m29b66_1 & x_m29b66_2;
   PP_m29_66X2Y1_Tbl: SmallMultTableP3x3r6XuYu_comb_uid68
      port map ( X => Y1X2_66_m29,
                 Y => PP66X2Y1_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w50_2 <= PP66X2Y1_m29(0); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w51_3 <= PP66X2Y1_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w52_3 <= PP66X2Y1_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w53_1 <= PP66X2Y1_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w54_2 <= PP66X2Y1_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w55_2 <= PP66X2Y1_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y1X3_66_m29 <= y_m29b66_1 & x_m29b66_3;
   PP_m29_66X3Y1_Tbl: SmallMultTableP3x3r6XuYu_comb_uid68
      port map ( X => Y1X3_66_m29,
                 Y => PP66X3Y1_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w53_2 <= PP66X3Y1_m29(0); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w54_3 <= PP66X3Y1_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w55_3 <= PP66X3Y1_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w56_1 <= PP66X3Y1_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w57_2 <= PP66X3Y1_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w58_2 <= PP66X3Y1_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y1X4_66_m29 <= y_m29b66_1 & x_m29b66_4;
   PP_m29_66X4Y1_Tbl: SmallMultTableP3x3r6XuYu_comb_uid68
      port map ( X => Y1X4_66_m29,
                 Y => PP66X4Y1_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w56_2 <= PP66X4Y1_m29(0); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w57_3 <= PP66X4Y1_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w58_3 <= PP66X4Y1_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w59_1 <= PP66X4Y1_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w60_2 <= PP66X4Y1_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w61_2 <= PP66X4Y1_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y1X5_66_m29 <= y_m29b66_1 & x_m29b66_5;
   PP_m29_66X5Y1_Tbl: SmallMultTableP3x3r6XuYu_comb_uid68
      port map ( X => Y1X5_66_m29,
                 Y => PP66X5Y1_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w59_2 <= PP66X5Y1_m29(0); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w60_3 <= PP66X5Y1_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w61_3 <= PP66X5Y1_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w62_1 <= PP66X5Y1_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w63_2 <= PP66X5Y1_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w64_2 <= PP66X5Y1_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y1X6_66_m29 <= y_m29b66_1 & x_m29b66_6;
   PP_m29_66X6Y1_Tbl: SmallMultTableP3x3r6XuYu_comb_uid68
      port map ( X => Y1X6_66_m29,
                 Y => PP66X6Y1_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w62_2 <= PP66X6Y1_m29(0); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w63_3 <= PP66X6Y1_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w64_3 <= PP66X6Y1_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w65_1 <= PP66X6Y1_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w66_2 <= PP66X6Y1_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w67_2 <= PP66X6Y1_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y1X7_66_m29 <= y_m29b66_1 & x_m29b66_7;
   PP_m29_66X7Y1_Tbl: SmallMultTableP3x3r6XuYu_comb_uid68
      port map ( X => Y1X7_66_m29,
                 Y => PP66X7Y1_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w65_2 <= PP66X7Y1_m29(0); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w66_3 <= PP66X7Y1_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w67_3 <= PP66X7Y1_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w68_2 <= PP66X7Y1_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w69_3 <= PP66X7Y1_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w70_3 <= PP66X7Y1_m29(5); -- cycle= 0 cp= 5.9176e-10

   -- code generated by IntMultiplier::buildHeapLogicOnly()
   -- buildheaplogiconly called for lsbX=18 lsbY=0 msbX=42 msbY=5
   Xp_m29b101 <= XX_m29(41 downto 18) & "";
   Yp_m29b101 <= YY_m29(4 downto 0) & "0";
   x_m29b101_0 <= Xp_m29b101(2 downto 0);
   x_m29b101_1 <= Xp_m29b101(5 downto 3);
   x_m29b101_2 <= Xp_m29b101(8 downto 6);
   x_m29b101_3 <= Xp_m29b101(11 downto 9);
   x_m29b101_4 <= Xp_m29b101(14 downto 12);
   x_m29b101_5 <= Xp_m29b101(17 downto 15);
   x_m29b101_6 <= Xp_m29b101(20 downto 18);
   x_m29b101_7 <= Xp_m29b101(23 downto 21);
   y_m29b101_0 <= Yp_m29b101(2 downto 0);
   y_m29b101_1 <= Yp_m29b101(5 downto 3);
   -- Partial product row number 0
   Y0X0_101_m29 <= y_m29b101_0 & x_m29b101_0;
   PP_m29_101X0Y0_Tbl: SmallMultTableP3x3r6XuYu_comb_uid103
      port map ( X => Y0X0_101_m29,
                 Y => PP101X0Y0_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w18_0 <= PP101X0Y0_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w19_0 <= PP101X0Y0_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w20_0 <= PP101X0Y0_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w21_0 <= PP101X0Y0_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w22_0 <= PP101X0Y0_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y0X1_101_m29 <= y_m29b101_0 & x_m29b101_1;
   PP_m29_101X1Y0_Tbl: SmallMultTableP3x3r6XuYu_comb_uid103
      port map ( X => Y0X1_101_m29,
                 Y => PP101X1Y0_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w21_1 <= PP101X1Y0_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w22_1 <= PP101X1Y0_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w23_0 <= PP101X1Y0_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w24_0 <= PP101X1Y0_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w25_0 <= PP101X1Y0_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y0X2_101_m29 <= y_m29b101_0 & x_m29b101_2;
   PP_m29_101X2Y0_Tbl: SmallMultTableP3x3r6XuYu_comb_uid103
      port map ( X => Y0X2_101_m29,
                 Y => PP101X2Y0_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w24_1 <= PP101X2Y0_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w25_1 <= PP101X2Y0_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w26_0 <= PP101X2Y0_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w27_0 <= PP101X2Y0_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w28_0 <= PP101X2Y0_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y0X3_101_m29 <= y_m29b101_0 & x_m29b101_3;
   PP_m29_101X3Y0_Tbl: SmallMultTableP3x3r6XuYu_comb_uid103
      port map ( X => Y0X3_101_m29,
                 Y => PP101X3Y0_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w27_1 <= PP101X3Y0_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w28_1 <= PP101X3Y0_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w29_0 <= PP101X3Y0_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w30_0 <= PP101X3Y0_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w31_0 <= PP101X3Y0_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y0X4_101_m29 <= y_m29b101_0 & x_m29b101_4;
   PP_m29_101X4Y0_Tbl: SmallMultTableP3x3r6XuYu_comb_uid103
      port map ( X => Y0X4_101_m29,
                 Y => PP101X4Y0_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w30_1 <= PP101X4Y0_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w31_1 <= PP101X4Y0_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w32_0 <= PP101X4Y0_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w33_0 <= PP101X4Y0_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w34_0 <= PP101X4Y0_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y0X5_101_m29 <= y_m29b101_0 & x_m29b101_5;
   PP_m29_101X5Y0_Tbl: SmallMultTableP3x3r6XuYu_comb_uid103
      port map ( X => Y0X5_101_m29,
                 Y => PP101X5Y0_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w33_1 <= PP101X5Y0_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w34_1 <= PP101X5Y0_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w35_0 <= PP101X5Y0_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w36_0 <= PP101X5Y0_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w37_0 <= PP101X5Y0_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y0X6_101_m29 <= y_m29b101_0 & x_m29b101_6;
   PP_m29_101X6Y0_Tbl: SmallMultTableP3x3r6XuYu_comb_uid103
      port map ( X => Y0X6_101_m29,
                 Y => PP101X6Y0_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w36_1 <= PP101X6Y0_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w37_1 <= PP101X6Y0_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w38_0 <= PP101X6Y0_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w39_0 <= PP101X6Y0_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w40_0 <= PP101X6Y0_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y0X7_101_m29 <= y_m29b101_0 & x_m29b101_7;
   PP_m29_101X7Y0_Tbl: SmallMultTableP3x3r6XuYu_comb_uid103
      port map ( X => Y0X7_101_m29,
                 Y => PP101X7Y0_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w39_1 <= PP101X7Y0_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w40_1 <= PP101X7Y0_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w41_0 <= PP101X7Y0_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w42_1 <= PP101X7Y0_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w43_1 <= PP101X7Y0_m29(5); -- cycle= 0 cp= 5.9176e-10

   -- Partial product row number 1
   Y1X0_101_m29 <= y_m29b101_1 & x_m29b101_0;
   PP_m29_101X0Y1_Tbl: SmallMultTableP3x3r6XuYu_comb_uid103
      port map ( X => Y1X0_101_m29,
                 Y => PP101X0Y1_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w20_1 <= PP101X0Y1_m29(0); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w21_2 <= PP101X0Y1_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w22_2 <= PP101X0Y1_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w23_1 <= PP101X0Y1_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w24_2 <= PP101X0Y1_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w25_2 <= PP101X0Y1_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y1X1_101_m29 <= y_m29b101_1 & x_m29b101_1;
   PP_m29_101X1Y1_Tbl: SmallMultTableP3x3r6XuYu_comb_uid103
      port map ( X => Y1X1_101_m29,
                 Y => PP101X1Y1_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w23_2 <= PP101X1Y1_m29(0); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w24_3 <= PP101X1Y1_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w25_3 <= PP101X1Y1_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w26_1 <= PP101X1Y1_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w27_2 <= PP101X1Y1_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w28_2 <= PP101X1Y1_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y1X2_101_m29 <= y_m29b101_1 & x_m29b101_2;
   PP_m29_101X2Y1_Tbl: SmallMultTableP3x3r6XuYu_comb_uid103
      port map ( X => Y1X2_101_m29,
                 Y => PP101X2Y1_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w26_2 <= PP101X2Y1_m29(0); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w27_3 <= PP101X2Y1_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w28_3 <= PP101X2Y1_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w29_1 <= PP101X2Y1_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w30_2 <= PP101X2Y1_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w31_2 <= PP101X2Y1_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y1X3_101_m29 <= y_m29b101_1 & x_m29b101_3;
   PP_m29_101X3Y1_Tbl: SmallMultTableP3x3r6XuYu_comb_uid103
      port map ( X => Y1X3_101_m29,
                 Y => PP101X3Y1_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w29_2 <= PP101X3Y1_m29(0); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w30_3 <= PP101X3Y1_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w31_3 <= PP101X3Y1_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w32_1 <= PP101X3Y1_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w33_2 <= PP101X3Y1_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w34_2 <= PP101X3Y1_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y1X4_101_m29 <= y_m29b101_1 & x_m29b101_4;
   PP_m29_101X4Y1_Tbl: SmallMultTableP3x3r6XuYu_comb_uid103
      port map ( X => Y1X4_101_m29,
                 Y => PP101X4Y1_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w32_2 <= PP101X4Y1_m29(0); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w33_3 <= PP101X4Y1_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w34_3 <= PP101X4Y1_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w35_1 <= PP101X4Y1_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w36_2 <= PP101X4Y1_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w37_2 <= PP101X4Y1_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y1X5_101_m29 <= y_m29b101_1 & x_m29b101_5;
   PP_m29_101X5Y1_Tbl: SmallMultTableP3x3r6XuYu_comb_uid103
      port map ( X => Y1X5_101_m29,
                 Y => PP101X5Y1_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w35_2 <= PP101X5Y1_m29(0); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w36_3 <= PP101X5Y1_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w37_3 <= PP101X5Y1_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w38_1 <= PP101X5Y1_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w39_2 <= PP101X5Y1_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w40_2 <= PP101X5Y1_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y1X6_101_m29 <= y_m29b101_1 & x_m29b101_6;
   PP_m29_101X6Y1_Tbl: SmallMultTableP3x3r6XuYu_comb_uid103
      port map ( X => Y1X6_101_m29,
                 Y => PP101X6Y1_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w38_2 <= PP101X6Y1_m29(0); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w39_3 <= PP101X6Y1_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w40_3 <= PP101X6Y1_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w41_1 <= PP101X6Y1_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w42_2 <= PP101X6Y1_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w43_2 <= PP101X6Y1_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y1X7_101_m29 <= y_m29b101_1 & x_m29b101_7;
   PP_m29_101X7Y1_Tbl: SmallMultTableP3x3r6XuYu_comb_uid103
      port map ( X => Y1X7_101_m29,
                 Y => PP101X7Y1_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w41_2 <= PP101X7Y1_m29(0); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w42_3 <= PP101X7Y1_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w43_3 <= PP101X7Y1_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w44_2 <= PP101X7Y1_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w45_3 <= PP101X7Y1_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w46_3 <= PP101X7Y1_m29(5); -- cycle= 0 cp= 5.9176e-10

   -- code generated by IntMultiplier::buildHeapLogicOnly()
   -- buildheaplogiconly called for lsbX=0 lsbY=0 msbX=18 msbY=5
   Xp_m29b136 <= XX_m29(17 downto 0) & "";
   Yp_m29b136 <= YY_m29(4 downto 0) & "0";
   x_m29b136_0 <= Xp_m29b136(2 downto 0);
   x_m29b136_1 <= Xp_m29b136(5 downto 3);
   x_m29b136_2 <= Xp_m29b136(8 downto 6);
   x_m29b136_3 <= Xp_m29b136(11 downto 9);
   x_m29b136_4 <= Xp_m29b136(14 downto 12);
   x_m29b136_5 <= Xp_m29b136(17 downto 15);
   y_m29b136_0 <= Yp_m29b136(2 downto 0);
   y_m29b136_1 <= Yp_m29b136(5 downto 3);
   -- Partial product row number 0
   Y0X0_136_m29 <= y_m29b136_0 & x_m29b136_0;
   PP_m29_136X0Y0_Tbl: SmallMultTableP3x3r6XuYu_comb_uid138
      port map ( X => Y0X0_136_m29,
                 Y => PP136X0Y0_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w0_0 <= PP136X0Y0_m29(1); -- cycle= 0 cp= 5.7432e-10
   heap_bh30_w1_0 <= PP136X0Y0_m29(2); -- cycle= 0 cp= 5.7432e-10
   heap_bh30_w2_0 <= PP136X0Y0_m29(3); -- cycle= 0 cp= 5.7432e-10
   heap_bh30_w3_0 <= PP136X0Y0_m29(4); -- cycle= 0 cp= 5.7432e-10
   heap_bh30_w4_0 <= PP136X0Y0_m29(5); -- cycle= 0 cp= 5.7432e-10

   Y0X1_136_m29 <= y_m29b136_0 & x_m29b136_1;
   PP_m29_136X1Y0_Tbl: SmallMultTableP3x3r6XuYu_comb_uid138
      port map ( X => Y0X1_136_m29,
                 Y => PP136X1Y0_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w3_1 <= PP136X1Y0_m29(1); -- cycle= 0 cp= 5.7432e-10
   heap_bh30_w4_1 <= PP136X1Y0_m29(2); -- cycle= 0 cp= 5.7432e-10
   heap_bh30_w5_0 <= PP136X1Y0_m29(3); -- cycle= 0 cp= 5.7432e-10
   heap_bh30_w6_0 <= PP136X1Y0_m29(4); -- cycle= 0 cp= 5.7432e-10
   heap_bh30_w7_0 <= PP136X1Y0_m29(5); -- cycle= 0 cp= 5.7432e-10

   Y0X2_136_m29 <= y_m29b136_0 & x_m29b136_2;
   PP_m29_136X2Y0_Tbl: SmallMultTableP3x3r6XuYu_comb_uid138
      port map ( X => Y0X2_136_m29,
                 Y => PP136X2Y0_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w6_1 <= PP136X2Y0_m29(1); -- cycle= 0 cp= 5.7432e-10
   heap_bh30_w7_1 <= PP136X2Y0_m29(2); -- cycle= 0 cp= 5.7432e-10
   heap_bh30_w8_0 <= PP136X2Y0_m29(3); -- cycle= 0 cp= 5.7432e-10
   heap_bh30_w9_0 <= PP136X2Y0_m29(4); -- cycle= 0 cp= 5.7432e-10
   heap_bh30_w10_0 <= PP136X2Y0_m29(5); -- cycle= 0 cp= 5.7432e-10

   Y0X3_136_m29 <= y_m29b136_0 & x_m29b136_3;
   PP_m29_136X3Y0_Tbl: SmallMultTableP3x3r6XuYu_comb_uid138
      port map ( X => Y0X3_136_m29,
                 Y => PP136X3Y0_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w9_1 <= PP136X3Y0_m29(1); -- cycle= 0 cp= 5.7432e-10
   heap_bh30_w10_1 <= PP136X3Y0_m29(2); -- cycle= 0 cp= 5.7432e-10
   heap_bh30_w11_0 <= PP136X3Y0_m29(3); -- cycle= 0 cp= 5.7432e-10
   heap_bh30_w12_0 <= PP136X3Y0_m29(4); -- cycle= 0 cp= 5.7432e-10
   heap_bh30_w13_0 <= PP136X3Y0_m29(5); -- cycle= 0 cp= 5.7432e-10

   Y0X4_136_m29 <= y_m29b136_0 & x_m29b136_4;
   PP_m29_136X4Y0_Tbl: SmallMultTableP3x3r6XuYu_comb_uid138
      port map ( X => Y0X4_136_m29,
                 Y => PP136X4Y0_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w12_1 <= PP136X4Y0_m29(1); -- cycle= 0 cp= 5.7432e-10
   heap_bh30_w13_1 <= PP136X4Y0_m29(2); -- cycle= 0 cp= 5.7432e-10
   heap_bh30_w14_0 <= PP136X4Y0_m29(3); -- cycle= 0 cp= 5.7432e-10
   heap_bh30_w15_0 <= PP136X4Y0_m29(4); -- cycle= 0 cp= 5.7432e-10
   heap_bh30_w16_0 <= PP136X4Y0_m29(5); -- cycle= 0 cp= 5.7432e-10

   Y0X5_136_m29 <= y_m29b136_0 & x_m29b136_5;
   PP_m29_136X5Y0_Tbl: SmallMultTableP3x3r6XuYu_comb_uid138
      port map ( X => Y0X5_136_m29,
                 Y => PP136X5Y0_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w15_1 <= PP136X5Y0_m29(1); -- cycle= 0 cp= 5.7432e-10
   heap_bh30_w16_1 <= PP136X5Y0_m29(2); -- cycle= 0 cp= 5.7432e-10
   heap_bh30_w17_0 <= PP136X5Y0_m29(3); -- cycle= 0 cp= 5.7432e-10
   heap_bh30_w18_1 <= PP136X5Y0_m29(4); -- cycle= 0 cp= 5.7432e-10
   heap_bh30_w19_1 <= PP136X5Y0_m29(5); -- cycle= 0 cp= 5.7432e-10

   -- Partial product row number 1
   Y1X0_136_m29 <= y_m29b136_1 & x_m29b136_0;
   PP_m29_136X0Y1_Tbl: SmallMultTableP3x3r6XuYu_comb_uid138
      port map ( X => Y1X0_136_m29,
                 Y => PP136X0Y1_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w2_1 <= PP136X0Y1_m29(0); -- cycle= 0 cp= 5.7432e-10
   heap_bh30_w3_2 <= PP136X0Y1_m29(1); -- cycle= 0 cp= 5.7432e-10
   heap_bh30_w4_2 <= PP136X0Y1_m29(2); -- cycle= 0 cp= 5.7432e-10
   heap_bh30_w5_1 <= PP136X0Y1_m29(3); -- cycle= 0 cp= 5.7432e-10
   heap_bh30_w6_2 <= PP136X0Y1_m29(4); -- cycle= 0 cp= 5.7432e-10
   heap_bh30_w7_2 <= PP136X0Y1_m29(5); -- cycle= 0 cp= 5.7432e-10

   Y1X1_136_m29 <= y_m29b136_1 & x_m29b136_1;
   PP_m29_136X1Y1_Tbl: SmallMultTableP3x3r6XuYu_comb_uid138
      port map ( X => Y1X1_136_m29,
                 Y => PP136X1Y1_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w5_2 <= PP136X1Y1_m29(0); -- cycle= 0 cp= 5.7432e-10
   heap_bh30_w6_3 <= PP136X1Y1_m29(1); -- cycle= 0 cp= 5.7432e-10
   heap_bh30_w7_3 <= PP136X1Y1_m29(2); -- cycle= 0 cp= 5.7432e-10
   heap_bh30_w8_1 <= PP136X1Y1_m29(3); -- cycle= 0 cp= 5.7432e-10
   heap_bh30_w9_2 <= PP136X1Y1_m29(4); -- cycle= 0 cp= 5.7432e-10
   heap_bh30_w10_2 <= PP136X1Y1_m29(5); -- cycle= 0 cp= 5.7432e-10

   Y1X2_136_m29 <= y_m29b136_1 & x_m29b136_2;
   PP_m29_136X2Y1_Tbl: SmallMultTableP3x3r6XuYu_comb_uid138
      port map ( X => Y1X2_136_m29,
                 Y => PP136X2Y1_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w8_2 <= PP136X2Y1_m29(0); -- cycle= 0 cp= 5.7432e-10
   heap_bh30_w9_3 <= PP136X2Y1_m29(1); -- cycle= 0 cp= 5.7432e-10
   heap_bh30_w10_3 <= PP136X2Y1_m29(2); -- cycle= 0 cp= 5.7432e-10
   heap_bh30_w11_1 <= PP136X2Y1_m29(3); -- cycle= 0 cp= 5.7432e-10
   heap_bh30_w12_2 <= PP136X2Y1_m29(4); -- cycle= 0 cp= 5.7432e-10
   heap_bh30_w13_2 <= PP136X2Y1_m29(5); -- cycle= 0 cp= 5.7432e-10

   Y1X3_136_m29 <= y_m29b136_1 & x_m29b136_3;
   PP_m29_136X3Y1_Tbl: SmallMultTableP3x3r6XuYu_comb_uid138
      port map ( X => Y1X3_136_m29,
                 Y => PP136X3Y1_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w11_2 <= PP136X3Y1_m29(0); -- cycle= 0 cp= 5.7432e-10
   heap_bh30_w12_3 <= PP136X3Y1_m29(1); -- cycle= 0 cp= 5.7432e-10
   heap_bh30_w13_3 <= PP136X3Y1_m29(2); -- cycle= 0 cp= 5.7432e-10
   heap_bh30_w14_1 <= PP136X3Y1_m29(3); -- cycle= 0 cp= 5.7432e-10
   heap_bh30_w15_2 <= PP136X3Y1_m29(4); -- cycle= 0 cp= 5.7432e-10
   heap_bh30_w16_2 <= PP136X3Y1_m29(5); -- cycle= 0 cp= 5.7432e-10

   Y1X4_136_m29 <= y_m29b136_1 & x_m29b136_4;
   PP_m29_136X4Y1_Tbl: SmallMultTableP3x3r6XuYu_comb_uid138
      port map ( X => Y1X4_136_m29,
                 Y => PP136X4Y1_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w14_2 <= PP136X4Y1_m29(0); -- cycle= 0 cp= 5.7432e-10
   heap_bh30_w15_3 <= PP136X4Y1_m29(1); -- cycle= 0 cp= 5.7432e-10
   heap_bh30_w16_3 <= PP136X4Y1_m29(2); -- cycle= 0 cp= 5.7432e-10
   heap_bh30_w17_1 <= PP136X4Y1_m29(3); -- cycle= 0 cp= 5.7432e-10
   heap_bh30_w18_2 <= PP136X4Y1_m29(4); -- cycle= 0 cp= 5.7432e-10
   heap_bh30_w19_2 <= PP136X4Y1_m29(5); -- cycle= 0 cp= 5.7432e-10

   Y1X5_136_m29 <= y_m29b136_1 & x_m29b136_5;
   PP_m29_136X5Y1_Tbl: SmallMultTableP3x3r6XuYu_comb_uid138
      port map ( X => Y1X5_136_m29,
                 Y => PP136X5Y1_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w17_2 <= PP136X5Y1_m29(0); -- cycle= 0 cp= 5.7432e-10
   heap_bh30_w18_3 <= PP136X5Y1_m29(1); -- cycle= 0 cp= 5.7432e-10
   heap_bh30_w19_3 <= PP136X5Y1_m29(2); -- cycle= 0 cp= 5.7432e-10
   heap_bh30_w20_2 <= PP136X5Y1_m29(3); -- cycle= 0 cp= 5.7432e-10
   heap_bh30_w21_3 <= PP136X5Y1_m29(4); -- cycle= 0 cp= 5.7432e-10
   heap_bh30_w22_3 <= PP136X5Y1_m29(5); -- cycle= 0 cp= 5.7432e-10

   
   -- Beginning of code generated by BitHeap::generateCompressorVHDL
   -- code generated by BitHeap::generateSupertileVHDL()
   DSP_bh30_ch0_0 <= std_logic_vector(unsigned("" & XX_m29(89 downto 66) & "") * unsigned("" & YY_m29(89 downto 73) & ""));
   heap_bh30_w179_0 <= DSP_bh30_ch0_0(40); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w178_0 <= DSP_bh30_ch0_0(39); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w177_0 <= DSP_bh30_ch0_0(38); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w176_0 <= DSP_bh30_ch0_0(37); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w175_0 <= DSP_bh30_ch0_0(36); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w174_0 <= DSP_bh30_ch0_0(35); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w173_0 <= DSP_bh30_ch0_0(34); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w172_0 <= DSP_bh30_ch0_0(33); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w171_0 <= DSP_bh30_ch0_0(32); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w170_0 <= DSP_bh30_ch0_0(31); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w169_0 <= DSP_bh30_ch0_0(30); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w168_0 <= DSP_bh30_ch0_0(29); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w167_0 <= DSP_bh30_ch0_0(28); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w166_0 <= DSP_bh30_ch0_0(27); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w165_0 <= DSP_bh30_ch0_0(26); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w164_0 <= DSP_bh30_ch0_0(25); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w163_0 <= DSP_bh30_ch0_0(24); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w162_0 <= DSP_bh30_ch0_0(23); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w161_0 <= DSP_bh30_ch0_0(22); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w160_0 <= DSP_bh30_ch0_0(21); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w159_0 <= DSP_bh30_ch0_0(20); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w158_0 <= DSP_bh30_ch0_0(19); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w157_0 <= DSP_bh30_ch0_0(18); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w156_0 <= DSP_bh30_ch0_0(17); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w155_0 <= DSP_bh30_ch0_0(16); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w154_0 <= DSP_bh30_ch0_0(15); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w153_0 <= DSP_bh30_ch0_0(14); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w152_0 <= DSP_bh30_ch0_0(13); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w151_0 <= DSP_bh30_ch0_0(12); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w150_0 <= DSP_bh30_ch0_0(11); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w149_0 <= DSP_bh30_ch0_0(10); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w148_0 <= DSP_bh30_ch0_0(9); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w147_0 <= DSP_bh30_ch0_0(8); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w146_0 <= DSP_bh30_ch0_0(7); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w145_0 <= DSP_bh30_ch0_0(6); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w144_0 <= DSP_bh30_ch0_0(5); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w143_0 <= DSP_bh30_ch0_0(4); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w142_0 <= DSP_bh30_ch0_0(3); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w141_0 <= DSP_bh30_ch0_0(2); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w140_0 <= DSP_bh30_ch0_0(1); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w139_0 <= DSP_bh30_ch0_0(0); -- cycle= 0 cp= 2.387e-09
   DSP_bh30_ch1_0 <= std_logic_vector(unsigned("" & XX_m29(65 downto 42) & "") * unsigned("" & YY_m29(89 downto 73) & ""));
   heap_bh30_w155_1 <= DSP_bh30_ch1_0(40); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w154_1 <= DSP_bh30_ch1_0(39); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w153_1 <= DSP_bh30_ch1_0(38); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w152_1 <= DSP_bh30_ch1_0(37); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w151_1 <= DSP_bh30_ch1_0(36); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w150_1 <= DSP_bh30_ch1_0(35); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w149_1 <= DSP_bh30_ch1_0(34); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w148_1 <= DSP_bh30_ch1_0(33); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w147_1 <= DSP_bh30_ch1_0(32); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w146_1 <= DSP_bh30_ch1_0(31); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w145_1 <= DSP_bh30_ch1_0(30); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w144_1 <= DSP_bh30_ch1_0(29); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w143_1 <= DSP_bh30_ch1_0(28); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w142_1 <= DSP_bh30_ch1_0(27); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w141_1 <= DSP_bh30_ch1_0(26); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w140_1 <= DSP_bh30_ch1_0(25); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w139_1 <= DSP_bh30_ch1_0(24); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w138_0 <= DSP_bh30_ch1_0(23); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w137_0 <= DSP_bh30_ch1_0(22); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w136_0 <= DSP_bh30_ch1_0(21); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w135_0 <= DSP_bh30_ch1_0(20); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w134_0 <= DSP_bh30_ch1_0(19); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w133_0 <= DSP_bh30_ch1_0(18); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w132_0 <= DSP_bh30_ch1_0(17); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w131_0 <= DSP_bh30_ch1_0(16); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w130_0 <= DSP_bh30_ch1_0(15); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w129_0 <= DSP_bh30_ch1_0(14); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w128_0 <= DSP_bh30_ch1_0(13); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w127_0 <= DSP_bh30_ch1_0(12); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w126_0 <= DSP_bh30_ch1_0(11); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w125_0 <= DSP_bh30_ch1_0(10); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w124_0 <= DSP_bh30_ch1_0(9); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w123_0 <= DSP_bh30_ch1_0(8); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w122_0 <= DSP_bh30_ch1_0(7); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w121_0 <= DSP_bh30_ch1_0(6); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w120_0 <= DSP_bh30_ch1_0(5); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w119_0 <= DSP_bh30_ch1_0(4); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w118_0 <= DSP_bh30_ch1_0(3); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w117_0 <= DSP_bh30_ch1_0(2); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w116_0 <= DSP_bh30_ch1_0(1); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w115_0 <= DSP_bh30_ch1_0(0); -- cycle= 0 cp= 2.387e-09
   DSP_bh30_ch2_0 <= std_logic_vector(unsigned("" & XX_m29(41 downto 18) & "") * unsigned("" & YY_m29(89 downto 73) & ""));
   heap_bh30_w131_1 <= DSP_bh30_ch2_0(40); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w130_1 <= DSP_bh30_ch2_0(39); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w129_1 <= DSP_bh30_ch2_0(38); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w128_1 <= DSP_bh30_ch2_0(37); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w127_1 <= DSP_bh30_ch2_0(36); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w126_1 <= DSP_bh30_ch2_0(35); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w125_1 <= DSP_bh30_ch2_0(34); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w124_1 <= DSP_bh30_ch2_0(33); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w123_1 <= DSP_bh30_ch2_0(32); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w122_1 <= DSP_bh30_ch2_0(31); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w121_1 <= DSP_bh30_ch2_0(30); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w120_1 <= DSP_bh30_ch2_0(29); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w119_1 <= DSP_bh30_ch2_0(28); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w118_1 <= DSP_bh30_ch2_0(27); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w117_1 <= DSP_bh30_ch2_0(26); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w116_1 <= DSP_bh30_ch2_0(25); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w115_1 <= DSP_bh30_ch2_0(24); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w114_0 <= DSP_bh30_ch2_0(23); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w113_0 <= DSP_bh30_ch2_0(22); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w112_0 <= DSP_bh30_ch2_0(21); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w111_0 <= DSP_bh30_ch2_0(20); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w110_0 <= DSP_bh30_ch2_0(19); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w109_0 <= DSP_bh30_ch2_0(18); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w108_0 <= DSP_bh30_ch2_0(17); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w107_0 <= DSP_bh30_ch2_0(16); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w106_0 <= DSP_bh30_ch2_0(15); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w105_0 <= DSP_bh30_ch2_0(14); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w104_0 <= DSP_bh30_ch2_0(13); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w103_0 <= DSP_bh30_ch2_0(12); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w102_0 <= DSP_bh30_ch2_0(11); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w101_0 <= DSP_bh30_ch2_0(10); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w100_0 <= DSP_bh30_ch2_0(9); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w99_0 <= DSP_bh30_ch2_0(8); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w98_0 <= DSP_bh30_ch2_0(7); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w97_0 <= DSP_bh30_ch2_0(6); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w96_0 <= DSP_bh30_ch2_0(5); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w95_0 <= DSP_bh30_ch2_0(4); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w94_1 <= DSP_bh30_ch2_0(3); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w93_1 <= DSP_bh30_ch2_0(2); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w92_1 <= DSP_bh30_ch2_0(1); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w91_3 <= DSP_bh30_ch2_0(0); -- cycle= 0 cp= 2.387e-09
   DSP_bh30_ch3_0 <= std_logic_vector(unsigned("" & XX_m29(17 downto 0) & "000000") * unsigned("" & YY_m29(89 downto 73) & ""));
   heap_bh30_w107_1 <= DSP_bh30_ch3_0(40); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w106_1 <= DSP_bh30_ch3_0(39); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w105_1 <= DSP_bh30_ch3_0(38); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w104_1 <= DSP_bh30_ch3_0(37); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w103_1 <= DSP_bh30_ch3_0(36); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w102_1 <= DSP_bh30_ch3_0(35); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w101_1 <= DSP_bh30_ch3_0(34); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w100_1 <= DSP_bh30_ch3_0(33); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w99_1 <= DSP_bh30_ch3_0(32); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w98_1 <= DSP_bh30_ch3_0(31); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w97_1 <= DSP_bh30_ch3_0(30); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w96_1 <= DSP_bh30_ch3_0(29); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w95_1 <= DSP_bh30_ch3_0(28); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w94_2 <= DSP_bh30_ch3_0(27); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w93_2 <= DSP_bh30_ch3_0(26); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w92_2 <= DSP_bh30_ch3_0(25); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w91_4 <= DSP_bh30_ch3_0(24); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w90_3 <= DSP_bh30_ch3_0(23); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w89_3 <= DSP_bh30_ch3_0(22); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w88_4 <= DSP_bh30_ch3_0(21); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w87_4 <= DSP_bh30_ch3_0(20); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w86_3 <= DSP_bh30_ch3_0(19); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w85_4 <= DSP_bh30_ch3_0(18); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w84_4 <= DSP_bh30_ch3_0(17); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w83_3 <= DSP_bh30_ch3_0(16); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w82_4 <= DSP_bh30_ch3_0(15); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w81_4 <= DSP_bh30_ch3_0(14); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w80_3 <= DSP_bh30_ch3_0(13); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w79_4 <= DSP_bh30_ch3_0(12); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w78_4 <= DSP_bh30_ch3_0(11); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w77_3 <= DSP_bh30_ch3_0(10); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w76_4 <= DSP_bh30_ch3_0(9); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w75_4 <= DSP_bh30_ch3_0(8); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w74_3 <= DSP_bh30_ch3_0(7); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w73_4 <= DSP_bh30_ch3_0(6); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w72_4 <= DSP_bh30_ch3_0(5); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w71_3 <= DSP_bh30_ch3_0(4); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w70_4 <= DSP_bh30_ch3_0(3); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w69_4 <= DSP_bh30_ch3_0(2); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w68_3 <= DSP_bh30_ch3_0(1); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w67_4 <= DSP_bh30_ch3_0(0); -- cycle= 0 cp= 2.387e-09
   DSP_bh30_ch4_0 <= std_logic_vector(unsigned("" & XX_m29(89 downto 66) & "") * unsigned("" & YY_m29(72 downto 56) & ""));
   heap_bh30_w162_1 <= DSP_bh30_ch4_0(40); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w161_1 <= DSP_bh30_ch4_0(39); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w160_1 <= DSP_bh30_ch4_0(38); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w159_1 <= DSP_bh30_ch4_0(37); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w158_1 <= DSP_bh30_ch4_0(36); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w157_1 <= DSP_bh30_ch4_0(35); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w156_1 <= DSP_bh30_ch4_0(34); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w155_2 <= DSP_bh30_ch4_0(33); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w154_2 <= DSP_bh30_ch4_0(32); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w153_2 <= DSP_bh30_ch4_0(31); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w152_2 <= DSP_bh30_ch4_0(30); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w151_2 <= DSP_bh30_ch4_0(29); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w150_2 <= DSP_bh30_ch4_0(28); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w149_2 <= DSP_bh30_ch4_0(27); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w148_2 <= DSP_bh30_ch4_0(26); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w147_2 <= DSP_bh30_ch4_0(25); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w146_2 <= DSP_bh30_ch4_0(24); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w145_2 <= DSP_bh30_ch4_0(23); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w144_2 <= DSP_bh30_ch4_0(22); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w143_2 <= DSP_bh30_ch4_0(21); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w142_2 <= DSP_bh30_ch4_0(20); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w141_2 <= DSP_bh30_ch4_0(19); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w140_2 <= DSP_bh30_ch4_0(18); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w139_2 <= DSP_bh30_ch4_0(17); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w138_1 <= DSP_bh30_ch4_0(16); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w137_1 <= DSP_bh30_ch4_0(15); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w136_1 <= DSP_bh30_ch4_0(14); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w135_1 <= DSP_bh30_ch4_0(13); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w134_1 <= DSP_bh30_ch4_0(12); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w133_1 <= DSP_bh30_ch4_0(11); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w132_1 <= DSP_bh30_ch4_0(10); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w131_2 <= DSP_bh30_ch4_0(9); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w130_2 <= DSP_bh30_ch4_0(8); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w129_2 <= DSP_bh30_ch4_0(7); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w128_2 <= DSP_bh30_ch4_0(6); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w127_2 <= DSP_bh30_ch4_0(5); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w126_2 <= DSP_bh30_ch4_0(4); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w125_2 <= DSP_bh30_ch4_0(3); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w124_2 <= DSP_bh30_ch4_0(2); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w123_2 <= DSP_bh30_ch4_0(1); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w122_2 <= DSP_bh30_ch4_0(0); -- cycle= 0 cp= 2.387e-09
   DSP_bh30_ch5_0 <= std_logic_vector(unsigned("" & XX_m29(65 downto 42) & "") * unsigned("" & YY_m29(72 downto 56) & ""));
   heap_bh30_w138_2 <= DSP_bh30_ch5_0(40); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w137_2 <= DSP_bh30_ch5_0(39); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w136_2 <= DSP_bh30_ch5_0(38); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w135_2 <= DSP_bh30_ch5_0(37); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w134_2 <= DSP_bh30_ch5_0(36); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w133_2 <= DSP_bh30_ch5_0(35); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w132_2 <= DSP_bh30_ch5_0(34); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w131_3 <= DSP_bh30_ch5_0(33); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w130_3 <= DSP_bh30_ch5_0(32); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w129_3 <= DSP_bh30_ch5_0(31); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w128_3 <= DSP_bh30_ch5_0(30); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w127_3 <= DSP_bh30_ch5_0(29); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w126_3 <= DSP_bh30_ch5_0(28); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w125_3 <= DSP_bh30_ch5_0(27); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w124_3 <= DSP_bh30_ch5_0(26); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w123_3 <= DSP_bh30_ch5_0(25); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w122_3 <= DSP_bh30_ch5_0(24); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w121_2 <= DSP_bh30_ch5_0(23); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w120_2 <= DSP_bh30_ch5_0(22); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w119_2 <= DSP_bh30_ch5_0(21); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w118_2 <= DSP_bh30_ch5_0(20); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w117_2 <= DSP_bh30_ch5_0(19); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w116_2 <= DSP_bh30_ch5_0(18); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w115_2 <= DSP_bh30_ch5_0(17); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w114_1 <= DSP_bh30_ch5_0(16); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w113_1 <= DSP_bh30_ch5_0(15); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w112_1 <= DSP_bh30_ch5_0(14); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w111_1 <= DSP_bh30_ch5_0(13); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w110_1 <= DSP_bh30_ch5_0(12); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w109_1 <= DSP_bh30_ch5_0(11); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w108_1 <= DSP_bh30_ch5_0(10); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w107_2 <= DSP_bh30_ch5_0(9); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w106_2 <= DSP_bh30_ch5_0(8); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w105_2 <= DSP_bh30_ch5_0(7); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w104_2 <= DSP_bh30_ch5_0(6); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w103_2 <= DSP_bh30_ch5_0(5); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w102_2 <= DSP_bh30_ch5_0(4); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w101_2 <= DSP_bh30_ch5_0(3); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w100_2 <= DSP_bh30_ch5_0(2); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w99_2 <= DSP_bh30_ch5_0(1); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w98_2 <= DSP_bh30_ch5_0(0); -- cycle= 0 cp= 2.387e-09
   DSP_bh30_ch6_0 <= std_logic_vector(unsigned("" & XX_m29(41 downto 18) & "") * unsigned("" & YY_m29(72 downto 56) & ""));
   heap_bh30_w114_2 <= DSP_bh30_ch6_0(40); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w113_2 <= DSP_bh30_ch6_0(39); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w112_2 <= DSP_bh30_ch6_0(38); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w111_2 <= DSP_bh30_ch6_0(37); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w110_2 <= DSP_bh30_ch6_0(36); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w109_2 <= DSP_bh30_ch6_0(35); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w108_2 <= DSP_bh30_ch6_0(34); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w107_3 <= DSP_bh30_ch6_0(33); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w106_3 <= DSP_bh30_ch6_0(32); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w105_3 <= DSP_bh30_ch6_0(31); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w104_3 <= DSP_bh30_ch6_0(30); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w103_3 <= DSP_bh30_ch6_0(29); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w102_3 <= DSP_bh30_ch6_0(28); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w101_3 <= DSP_bh30_ch6_0(27); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w100_3 <= DSP_bh30_ch6_0(26); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w99_3 <= DSP_bh30_ch6_0(25); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w98_3 <= DSP_bh30_ch6_0(24); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w97_2 <= DSP_bh30_ch6_0(23); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w96_2 <= DSP_bh30_ch6_0(22); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w95_2 <= DSP_bh30_ch6_0(21); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w94_3 <= DSP_bh30_ch6_0(20); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w93_3 <= DSP_bh30_ch6_0(19); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w92_3 <= DSP_bh30_ch6_0(18); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w91_5 <= DSP_bh30_ch6_0(17); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w90_4 <= DSP_bh30_ch6_0(16); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w89_4 <= DSP_bh30_ch6_0(15); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w88_5 <= DSP_bh30_ch6_0(14); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w87_5 <= DSP_bh30_ch6_0(13); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w86_4 <= DSP_bh30_ch6_0(12); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w85_5 <= DSP_bh30_ch6_0(11); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w84_5 <= DSP_bh30_ch6_0(10); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w83_4 <= DSP_bh30_ch6_0(9); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w82_5 <= DSP_bh30_ch6_0(8); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w81_5 <= DSP_bh30_ch6_0(7); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w80_4 <= DSP_bh30_ch6_0(6); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w79_5 <= DSP_bh30_ch6_0(5); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w78_5 <= DSP_bh30_ch6_0(4); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w77_4 <= DSP_bh30_ch6_0(3); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w76_5 <= DSP_bh30_ch6_0(2); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w75_5 <= DSP_bh30_ch6_0(1); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w74_4 <= DSP_bh30_ch6_0(0); -- cycle= 0 cp= 2.387e-09
   DSP_bh30_ch7_0 <= std_logic_vector(unsigned("" & XX_m29(17 downto 0) & "000000") * unsigned("" & YY_m29(72 downto 56) & ""));
   heap_bh30_w90_5 <= DSP_bh30_ch7_0(40); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w89_5 <= DSP_bh30_ch7_0(39); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w88_6 <= DSP_bh30_ch7_0(38); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w87_6 <= DSP_bh30_ch7_0(37); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w86_5 <= DSP_bh30_ch7_0(36); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w85_6 <= DSP_bh30_ch7_0(35); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w84_6 <= DSP_bh30_ch7_0(34); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w83_5 <= DSP_bh30_ch7_0(33); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w82_6 <= DSP_bh30_ch7_0(32); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w81_6 <= DSP_bh30_ch7_0(31); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w80_5 <= DSP_bh30_ch7_0(30); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w79_6 <= DSP_bh30_ch7_0(29); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w78_6 <= DSP_bh30_ch7_0(28); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w77_5 <= DSP_bh30_ch7_0(27); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w76_6 <= DSP_bh30_ch7_0(26); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w75_6 <= DSP_bh30_ch7_0(25); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w74_5 <= DSP_bh30_ch7_0(24); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w73_5 <= DSP_bh30_ch7_0(23); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w72_5 <= DSP_bh30_ch7_0(22); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w71_4 <= DSP_bh30_ch7_0(21); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w70_5 <= DSP_bh30_ch7_0(20); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w69_5 <= DSP_bh30_ch7_0(19); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w68_4 <= DSP_bh30_ch7_0(18); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w67_5 <= DSP_bh30_ch7_0(17); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w66_4 <= DSP_bh30_ch7_0(16); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w65_3 <= DSP_bh30_ch7_0(15); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w64_4 <= DSP_bh30_ch7_0(14); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w63_4 <= DSP_bh30_ch7_0(13); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w62_3 <= DSP_bh30_ch7_0(12); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w61_4 <= DSP_bh30_ch7_0(11); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w60_4 <= DSP_bh30_ch7_0(10); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w59_3 <= DSP_bh30_ch7_0(9); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w58_4 <= DSP_bh30_ch7_0(8); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w57_4 <= DSP_bh30_ch7_0(7); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w56_3 <= DSP_bh30_ch7_0(6); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w55_4 <= DSP_bh30_ch7_0(5); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w54_4 <= DSP_bh30_ch7_0(4); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w53_3 <= DSP_bh30_ch7_0(3); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w52_4 <= DSP_bh30_ch7_0(2); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w51_4 <= DSP_bh30_ch7_0(1); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w50_3 <= DSP_bh30_ch7_0(0); -- cycle= 0 cp= 2.387e-09
   DSP_bh30_ch8_0 <= std_logic_vector(unsigned("" & XX_m29(89 downto 66) & "") * unsigned("" & YY_m29(55 downto 39) & ""));
   heap_bh30_w145_3 <= DSP_bh30_ch8_0(40); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w144_3 <= DSP_bh30_ch8_0(39); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w143_3 <= DSP_bh30_ch8_0(38); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w142_3 <= DSP_bh30_ch8_0(37); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w141_3 <= DSP_bh30_ch8_0(36); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w140_3 <= DSP_bh30_ch8_0(35); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w139_3 <= DSP_bh30_ch8_0(34); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w138_3 <= DSP_bh30_ch8_0(33); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w137_3 <= DSP_bh30_ch8_0(32); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w136_3 <= DSP_bh30_ch8_0(31); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w135_3 <= DSP_bh30_ch8_0(30); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w134_3 <= DSP_bh30_ch8_0(29); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w133_3 <= DSP_bh30_ch8_0(28); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w132_3 <= DSP_bh30_ch8_0(27); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w131_4 <= DSP_bh30_ch8_0(26); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w130_4 <= DSP_bh30_ch8_0(25); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w129_4 <= DSP_bh30_ch8_0(24); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w128_4 <= DSP_bh30_ch8_0(23); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w127_4 <= DSP_bh30_ch8_0(22); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w126_4 <= DSP_bh30_ch8_0(21); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w125_4 <= DSP_bh30_ch8_0(20); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w124_4 <= DSP_bh30_ch8_0(19); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w123_4 <= DSP_bh30_ch8_0(18); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w122_4 <= DSP_bh30_ch8_0(17); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w121_3 <= DSP_bh30_ch8_0(16); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w120_3 <= DSP_bh30_ch8_0(15); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w119_3 <= DSP_bh30_ch8_0(14); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w118_3 <= DSP_bh30_ch8_0(13); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w117_3 <= DSP_bh30_ch8_0(12); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w116_3 <= DSP_bh30_ch8_0(11); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w115_3 <= DSP_bh30_ch8_0(10); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w114_3 <= DSP_bh30_ch8_0(9); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w113_3 <= DSP_bh30_ch8_0(8); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w112_3 <= DSP_bh30_ch8_0(7); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w111_3 <= DSP_bh30_ch8_0(6); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w110_3 <= DSP_bh30_ch8_0(5); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w109_3 <= DSP_bh30_ch8_0(4); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w108_3 <= DSP_bh30_ch8_0(3); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w107_4 <= DSP_bh30_ch8_0(2); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w106_4 <= DSP_bh30_ch8_0(1); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w105_4 <= DSP_bh30_ch8_0(0); -- cycle= 0 cp= 2.387e-09
   DSP_bh30_ch9_0 <= std_logic_vector(unsigned("" & XX_m29(65 downto 42) & "") * unsigned("" & YY_m29(55 downto 39) & ""));
   heap_bh30_w121_4 <= DSP_bh30_ch9_0(40); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w120_4 <= DSP_bh30_ch9_0(39); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w119_4 <= DSP_bh30_ch9_0(38); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w118_4 <= DSP_bh30_ch9_0(37); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w117_4 <= DSP_bh30_ch9_0(36); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w116_4 <= DSP_bh30_ch9_0(35); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w115_4 <= DSP_bh30_ch9_0(34); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w114_4 <= DSP_bh30_ch9_0(33); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w113_4 <= DSP_bh30_ch9_0(32); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w112_4 <= DSP_bh30_ch9_0(31); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w111_4 <= DSP_bh30_ch9_0(30); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w110_4 <= DSP_bh30_ch9_0(29); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w109_4 <= DSP_bh30_ch9_0(28); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w108_4 <= DSP_bh30_ch9_0(27); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w107_5 <= DSP_bh30_ch9_0(26); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w106_5 <= DSP_bh30_ch9_0(25); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w105_5 <= DSP_bh30_ch9_0(24); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w104_4 <= DSP_bh30_ch9_0(23); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w103_4 <= DSP_bh30_ch9_0(22); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w102_4 <= DSP_bh30_ch9_0(21); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w101_4 <= DSP_bh30_ch9_0(20); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w100_4 <= DSP_bh30_ch9_0(19); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w99_4 <= DSP_bh30_ch9_0(18); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w98_4 <= DSP_bh30_ch9_0(17); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w97_3 <= DSP_bh30_ch9_0(16); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w96_3 <= DSP_bh30_ch9_0(15); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w95_3 <= DSP_bh30_ch9_0(14); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w94_4 <= DSP_bh30_ch9_0(13); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w93_4 <= DSP_bh30_ch9_0(12); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w92_4 <= DSP_bh30_ch9_0(11); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w91_6 <= DSP_bh30_ch9_0(10); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w90_6 <= DSP_bh30_ch9_0(9); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w89_6 <= DSP_bh30_ch9_0(8); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w88_7 <= DSP_bh30_ch9_0(7); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w87_7 <= DSP_bh30_ch9_0(6); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w86_6 <= DSP_bh30_ch9_0(5); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w85_7 <= DSP_bh30_ch9_0(4); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w84_7 <= DSP_bh30_ch9_0(3); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w83_6 <= DSP_bh30_ch9_0(2); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w82_7 <= DSP_bh30_ch9_0(1); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w81_7 <= DSP_bh30_ch9_0(0); -- cycle= 0 cp= 2.387e-09
   DSP_bh30_ch10_0 <= std_logic_vector(unsigned("" & XX_m29(41 downto 18) & "") * unsigned("" & YY_m29(55 downto 39) & ""));
   heap_bh30_w97_4 <= DSP_bh30_ch10_0(40); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w96_4 <= DSP_bh30_ch10_0(39); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w95_4 <= DSP_bh30_ch10_0(38); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w94_5 <= DSP_bh30_ch10_0(37); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w93_5 <= DSP_bh30_ch10_0(36); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w92_5 <= DSP_bh30_ch10_0(35); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w91_7 <= DSP_bh30_ch10_0(34); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w90_7 <= DSP_bh30_ch10_0(33); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w89_7 <= DSP_bh30_ch10_0(32); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w88_8 <= DSP_bh30_ch10_0(31); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w87_8 <= DSP_bh30_ch10_0(30); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w86_7 <= DSP_bh30_ch10_0(29); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w85_8 <= DSP_bh30_ch10_0(28); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w84_8 <= DSP_bh30_ch10_0(27); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w83_7 <= DSP_bh30_ch10_0(26); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w82_8 <= DSP_bh30_ch10_0(25); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w81_8 <= DSP_bh30_ch10_0(24); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w80_6 <= DSP_bh30_ch10_0(23); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w79_7 <= DSP_bh30_ch10_0(22); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w78_7 <= DSP_bh30_ch10_0(21); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w77_6 <= DSP_bh30_ch10_0(20); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w76_7 <= DSP_bh30_ch10_0(19); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w75_7 <= DSP_bh30_ch10_0(18); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w74_6 <= DSP_bh30_ch10_0(17); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w73_6 <= DSP_bh30_ch10_0(16); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w72_6 <= DSP_bh30_ch10_0(15); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w71_5 <= DSP_bh30_ch10_0(14); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w70_6 <= DSP_bh30_ch10_0(13); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w69_6 <= DSP_bh30_ch10_0(12); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w68_5 <= DSP_bh30_ch10_0(11); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w67_6 <= DSP_bh30_ch10_0(10); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w66_5 <= DSP_bh30_ch10_0(9); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w65_4 <= DSP_bh30_ch10_0(8); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w64_5 <= DSP_bh30_ch10_0(7); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w63_5 <= DSP_bh30_ch10_0(6); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w62_4 <= DSP_bh30_ch10_0(5); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w61_5 <= DSP_bh30_ch10_0(4); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w60_5 <= DSP_bh30_ch10_0(3); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w59_4 <= DSP_bh30_ch10_0(2); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w58_5 <= DSP_bh30_ch10_0(1); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w57_5 <= DSP_bh30_ch10_0(0); -- cycle= 0 cp= 2.387e-09
   DSP_bh30_ch11_0 <= std_logic_vector(unsigned("" & XX_m29(17 downto 0) & "000000") * unsigned("" & YY_m29(55 downto 39) & ""));
   heap_bh30_w73_7 <= DSP_bh30_ch11_0(40); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w72_7 <= DSP_bh30_ch11_0(39); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w71_6 <= DSP_bh30_ch11_0(38); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w70_7 <= DSP_bh30_ch11_0(37); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w69_7 <= DSP_bh30_ch11_0(36); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w68_6 <= DSP_bh30_ch11_0(35); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w67_7 <= DSP_bh30_ch11_0(34); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w66_6 <= DSP_bh30_ch11_0(33); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w65_5 <= DSP_bh30_ch11_0(32); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w64_6 <= DSP_bh30_ch11_0(31); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w63_6 <= DSP_bh30_ch11_0(30); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w62_5 <= DSP_bh30_ch11_0(29); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w61_6 <= DSP_bh30_ch11_0(28); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w60_6 <= DSP_bh30_ch11_0(27); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w59_5 <= DSP_bh30_ch11_0(26); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w58_6 <= DSP_bh30_ch11_0(25); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w57_6 <= DSP_bh30_ch11_0(24); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w56_4 <= DSP_bh30_ch11_0(23); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w55_5 <= DSP_bh30_ch11_0(22); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w54_5 <= DSP_bh30_ch11_0(21); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w53_4 <= DSP_bh30_ch11_0(20); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w52_5 <= DSP_bh30_ch11_0(19); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w51_5 <= DSP_bh30_ch11_0(18); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w50_4 <= DSP_bh30_ch11_0(17); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w49_4 <= DSP_bh30_ch11_0(16); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w48_4 <= DSP_bh30_ch11_0(15); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w47_3 <= DSP_bh30_ch11_0(14); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w46_4 <= DSP_bh30_ch11_0(13); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w45_4 <= DSP_bh30_ch11_0(12); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w44_3 <= DSP_bh30_ch11_0(11); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w43_4 <= DSP_bh30_ch11_0(10); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w42_4 <= DSP_bh30_ch11_0(9); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w41_3 <= DSP_bh30_ch11_0(8); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w40_4 <= DSP_bh30_ch11_0(7); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w39_4 <= DSP_bh30_ch11_0(6); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w38_3 <= DSP_bh30_ch11_0(5); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w37_4 <= DSP_bh30_ch11_0(4); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w36_4 <= DSP_bh30_ch11_0(3); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w35_3 <= DSP_bh30_ch11_0(2); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w34_4 <= DSP_bh30_ch11_0(1); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w33_4 <= DSP_bh30_ch11_0(0); -- cycle= 0 cp= 2.387e-09
   DSP_bh30_ch12_0 <= std_logic_vector(unsigned("" & XX_m29(89 downto 66) & "") * unsigned("" & YY_m29(38 downto 22) & ""));
   heap_bh30_w128_5 <= DSP_bh30_ch12_0(40); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w127_5 <= DSP_bh30_ch12_0(39); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w126_5 <= DSP_bh30_ch12_0(38); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w125_5 <= DSP_bh30_ch12_0(37); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w124_5 <= DSP_bh30_ch12_0(36); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w123_5 <= DSP_bh30_ch12_0(35); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w122_5 <= DSP_bh30_ch12_0(34); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w121_5 <= DSP_bh30_ch12_0(33); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w120_5 <= DSP_bh30_ch12_0(32); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w119_5 <= DSP_bh30_ch12_0(31); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w118_5 <= DSP_bh30_ch12_0(30); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w117_5 <= DSP_bh30_ch12_0(29); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w116_5 <= DSP_bh30_ch12_0(28); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w115_5 <= DSP_bh30_ch12_0(27); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w114_5 <= DSP_bh30_ch12_0(26); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w113_5 <= DSP_bh30_ch12_0(25); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w112_5 <= DSP_bh30_ch12_0(24); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w111_5 <= DSP_bh30_ch12_0(23); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w110_5 <= DSP_bh30_ch12_0(22); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w109_5 <= DSP_bh30_ch12_0(21); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w108_5 <= DSP_bh30_ch12_0(20); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w107_6 <= DSP_bh30_ch12_0(19); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w106_6 <= DSP_bh30_ch12_0(18); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w105_6 <= DSP_bh30_ch12_0(17); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w104_5 <= DSP_bh30_ch12_0(16); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w103_5 <= DSP_bh30_ch12_0(15); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w102_5 <= DSP_bh30_ch12_0(14); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w101_5 <= DSP_bh30_ch12_0(13); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w100_5 <= DSP_bh30_ch12_0(12); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w99_5 <= DSP_bh30_ch12_0(11); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w98_5 <= DSP_bh30_ch12_0(10); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w97_5 <= DSP_bh30_ch12_0(9); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w96_5 <= DSP_bh30_ch12_0(8); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w95_5 <= DSP_bh30_ch12_0(7); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w94_6 <= DSP_bh30_ch12_0(6); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w93_6 <= DSP_bh30_ch12_0(5); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w92_6 <= DSP_bh30_ch12_0(4); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w91_8 <= DSP_bh30_ch12_0(3); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w90_8 <= DSP_bh30_ch12_0(2); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w89_8 <= DSP_bh30_ch12_0(1); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w88_9 <= DSP_bh30_ch12_0(0); -- cycle= 0 cp= 2.387e-09
   DSP_bh30_ch13_0 <= std_logic_vector(unsigned("" & XX_m29(65 downto 42) & "") * unsigned("" & YY_m29(38 downto 22) & ""));
   heap_bh30_w104_6 <= DSP_bh30_ch13_0(40); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w103_6 <= DSP_bh30_ch13_0(39); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w102_6 <= DSP_bh30_ch13_0(38); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w101_6 <= DSP_bh30_ch13_0(37); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w100_6 <= DSP_bh30_ch13_0(36); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w99_6 <= DSP_bh30_ch13_0(35); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w98_6 <= DSP_bh30_ch13_0(34); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w97_6 <= DSP_bh30_ch13_0(33); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w96_6 <= DSP_bh30_ch13_0(32); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w95_6 <= DSP_bh30_ch13_0(31); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w94_7 <= DSP_bh30_ch13_0(30); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w93_7 <= DSP_bh30_ch13_0(29); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w92_7 <= DSP_bh30_ch13_0(28); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w91_9 <= DSP_bh30_ch13_0(27); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w90_9 <= DSP_bh30_ch13_0(26); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w89_9 <= DSP_bh30_ch13_0(25); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w88_10 <= DSP_bh30_ch13_0(24); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w87_9 <= DSP_bh30_ch13_0(23); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w86_8 <= DSP_bh30_ch13_0(22); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w85_9 <= DSP_bh30_ch13_0(21); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w84_9 <= DSP_bh30_ch13_0(20); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w83_8 <= DSP_bh30_ch13_0(19); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w82_9 <= DSP_bh30_ch13_0(18); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w81_9 <= DSP_bh30_ch13_0(17); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w80_7 <= DSP_bh30_ch13_0(16); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w79_8 <= DSP_bh30_ch13_0(15); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w78_8 <= DSP_bh30_ch13_0(14); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w77_7 <= DSP_bh30_ch13_0(13); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w76_8 <= DSP_bh30_ch13_0(12); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w75_8 <= DSP_bh30_ch13_0(11); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w74_7 <= DSP_bh30_ch13_0(10); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w73_8 <= DSP_bh30_ch13_0(9); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w72_8 <= DSP_bh30_ch13_0(8); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w71_7 <= DSP_bh30_ch13_0(7); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w70_8 <= DSP_bh30_ch13_0(6); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w69_8 <= DSP_bh30_ch13_0(5); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w68_7 <= DSP_bh30_ch13_0(4); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w67_8 <= DSP_bh30_ch13_0(3); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w66_7 <= DSP_bh30_ch13_0(2); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w65_6 <= DSP_bh30_ch13_0(1); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w64_7 <= DSP_bh30_ch13_0(0); -- cycle= 0 cp= 2.387e-09
   DSP_bh30_ch14_0 <= std_logic_vector(unsigned("" & XX_m29(41 downto 18) & "") * unsigned("" & YY_m29(38 downto 22) & ""));
   heap_bh30_w80_8 <= DSP_bh30_ch14_0(40); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w79_9 <= DSP_bh30_ch14_0(39); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w78_9 <= DSP_bh30_ch14_0(38); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w77_8 <= DSP_bh30_ch14_0(37); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w76_9 <= DSP_bh30_ch14_0(36); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w75_9 <= DSP_bh30_ch14_0(35); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w74_8 <= DSP_bh30_ch14_0(34); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w73_9 <= DSP_bh30_ch14_0(33); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w72_9 <= DSP_bh30_ch14_0(32); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w71_8 <= DSP_bh30_ch14_0(31); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w70_9 <= DSP_bh30_ch14_0(30); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w69_9 <= DSP_bh30_ch14_0(29); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w68_8 <= DSP_bh30_ch14_0(28); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w67_9 <= DSP_bh30_ch14_0(27); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w66_8 <= DSP_bh30_ch14_0(26); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w65_7 <= DSP_bh30_ch14_0(25); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w64_8 <= DSP_bh30_ch14_0(24); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w63_7 <= DSP_bh30_ch14_0(23); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w62_6 <= DSP_bh30_ch14_0(22); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w61_7 <= DSP_bh30_ch14_0(21); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w60_7 <= DSP_bh30_ch14_0(20); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w59_6 <= DSP_bh30_ch14_0(19); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w58_7 <= DSP_bh30_ch14_0(18); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w57_7 <= DSP_bh30_ch14_0(17); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w56_5 <= DSP_bh30_ch14_0(16); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w55_6 <= DSP_bh30_ch14_0(15); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w54_6 <= DSP_bh30_ch14_0(14); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w53_5 <= DSP_bh30_ch14_0(13); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w52_6 <= DSP_bh30_ch14_0(12); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w51_6 <= DSP_bh30_ch14_0(11); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w50_5 <= DSP_bh30_ch14_0(10); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w49_5 <= DSP_bh30_ch14_0(9); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w48_5 <= DSP_bh30_ch14_0(8); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w47_4 <= DSP_bh30_ch14_0(7); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w46_5 <= DSP_bh30_ch14_0(6); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w45_5 <= DSP_bh30_ch14_0(5); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w44_4 <= DSP_bh30_ch14_0(4); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w43_5 <= DSP_bh30_ch14_0(3); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w42_5 <= DSP_bh30_ch14_0(2); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w41_4 <= DSP_bh30_ch14_0(1); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w40_5 <= DSP_bh30_ch14_0(0); -- cycle= 0 cp= 2.387e-09
   DSP_bh30_ch15_0 <= std_logic_vector(unsigned("" & XX_m29(17 downto 0) & "000000") * unsigned("" & YY_m29(38 downto 22) & ""));
   heap_bh30_w56_6 <= DSP_bh30_ch15_0(40); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w55_7 <= DSP_bh30_ch15_0(39); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w54_7 <= DSP_bh30_ch15_0(38); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w53_6 <= DSP_bh30_ch15_0(37); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w52_7 <= DSP_bh30_ch15_0(36); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w51_7 <= DSP_bh30_ch15_0(35); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w50_6 <= DSP_bh30_ch15_0(34); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w49_6 <= DSP_bh30_ch15_0(33); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w48_6 <= DSP_bh30_ch15_0(32); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w47_5 <= DSP_bh30_ch15_0(31); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w46_6 <= DSP_bh30_ch15_0(30); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w45_6 <= DSP_bh30_ch15_0(29); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w44_5 <= DSP_bh30_ch15_0(28); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w43_6 <= DSP_bh30_ch15_0(27); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w42_6 <= DSP_bh30_ch15_0(26); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w41_5 <= DSP_bh30_ch15_0(25); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w40_6 <= DSP_bh30_ch15_0(24); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w39_5 <= DSP_bh30_ch15_0(23); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w38_4 <= DSP_bh30_ch15_0(22); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w37_5 <= DSP_bh30_ch15_0(21); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w36_5 <= DSP_bh30_ch15_0(20); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w35_4 <= DSP_bh30_ch15_0(19); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w34_5 <= DSP_bh30_ch15_0(18); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w33_5 <= DSP_bh30_ch15_0(17); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w32_3 <= DSP_bh30_ch15_0(16); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w31_4 <= DSP_bh30_ch15_0(15); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w30_4 <= DSP_bh30_ch15_0(14); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w29_3 <= DSP_bh30_ch15_0(13); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w28_4 <= DSP_bh30_ch15_0(12); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w27_4 <= DSP_bh30_ch15_0(11); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w26_3 <= DSP_bh30_ch15_0(10); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w25_4 <= DSP_bh30_ch15_0(9); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w24_4 <= DSP_bh30_ch15_0(8); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w23_3 <= DSP_bh30_ch15_0(7); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w22_4 <= DSP_bh30_ch15_0(6); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w21_4 <= DSP_bh30_ch15_0(5); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w20_3 <= DSP_bh30_ch15_0(4); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w19_4 <= DSP_bh30_ch15_0(3); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w18_4 <= DSP_bh30_ch15_0(2); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w17_3 <= DSP_bh30_ch15_0(1); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w16_4 <= DSP_bh30_ch15_0(0); -- cycle= 0 cp= 2.387e-09
   DSP_bh30_ch16_0 <= std_logic_vector(unsigned("" & XX_m29(89 downto 66) & "") * unsigned("" & YY_m29(21 downto 5) & ""));
   heap_bh30_w111_6 <= DSP_bh30_ch16_0(40); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w110_6 <= DSP_bh30_ch16_0(39); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w109_6 <= DSP_bh30_ch16_0(38); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w108_6 <= DSP_bh30_ch16_0(37); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w107_7 <= DSP_bh30_ch16_0(36); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w106_7 <= DSP_bh30_ch16_0(35); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w105_7 <= DSP_bh30_ch16_0(34); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w104_7 <= DSP_bh30_ch16_0(33); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w103_7 <= DSP_bh30_ch16_0(32); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w102_7 <= DSP_bh30_ch16_0(31); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w101_7 <= DSP_bh30_ch16_0(30); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w100_7 <= DSP_bh30_ch16_0(29); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w99_7 <= DSP_bh30_ch16_0(28); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w98_7 <= DSP_bh30_ch16_0(27); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w97_7 <= DSP_bh30_ch16_0(26); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w96_7 <= DSP_bh30_ch16_0(25); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w95_7 <= DSP_bh30_ch16_0(24); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w94_8 <= DSP_bh30_ch16_0(23); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w93_8 <= DSP_bh30_ch16_0(22); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w92_8 <= DSP_bh30_ch16_0(21); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w91_10 <= DSP_bh30_ch16_0(20); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w90_10 <= DSP_bh30_ch16_0(19); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w89_10 <= DSP_bh30_ch16_0(18); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w88_11 <= DSP_bh30_ch16_0(17); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w87_10 <= DSP_bh30_ch16_0(16); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w86_9 <= DSP_bh30_ch16_0(15); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w85_10 <= DSP_bh30_ch16_0(14); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w84_10 <= DSP_bh30_ch16_0(13); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w83_9 <= DSP_bh30_ch16_0(12); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w82_10 <= DSP_bh30_ch16_0(11); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w81_10 <= DSP_bh30_ch16_0(10); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w80_9 <= DSP_bh30_ch16_0(9); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w79_10 <= DSP_bh30_ch16_0(8); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w78_10 <= DSP_bh30_ch16_0(7); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w77_9 <= DSP_bh30_ch16_0(6); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w76_10 <= DSP_bh30_ch16_0(5); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w75_10 <= DSP_bh30_ch16_0(4); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w74_9 <= DSP_bh30_ch16_0(3); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w73_10 <= DSP_bh30_ch16_0(2); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w72_10 <= DSP_bh30_ch16_0(1); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w71_9 <= DSP_bh30_ch16_0(0); -- cycle= 0 cp= 2.387e-09
   DSP_bh30_ch17_0 <= std_logic_vector(unsigned("" & XX_m29(65 downto 42) & "") * unsigned("" & YY_m29(21 downto 5) & ""));
   heap_bh30_w87_11 <= DSP_bh30_ch17_0(40); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w86_10 <= DSP_bh30_ch17_0(39); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w85_11 <= DSP_bh30_ch17_0(38); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w84_11 <= DSP_bh30_ch17_0(37); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w83_10 <= DSP_bh30_ch17_0(36); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w82_11 <= DSP_bh30_ch17_0(35); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w81_11 <= DSP_bh30_ch17_0(34); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w80_10 <= DSP_bh30_ch17_0(33); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w79_11 <= DSP_bh30_ch17_0(32); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w78_11 <= DSP_bh30_ch17_0(31); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w77_10 <= DSP_bh30_ch17_0(30); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w76_11 <= DSP_bh30_ch17_0(29); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w75_11 <= DSP_bh30_ch17_0(28); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w74_10 <= DSP_bh30_ch17_0(27); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w73_11 <= DSP_bh30_ch17_0(26); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w72_11 <= DSP_bh30_ch17_0(25); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w71_10 <= DSP_bh30_ch17_0(24); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w70_10 <= DSP_bh30_ch17_0(23); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w69_10 <= DSP_bh30_ch17_0(22); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w68_9 <= DSP_bh30_ch17_0(21); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w67_10 <= DSP_bh30_ch17_0(20); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w66_9 <= DSP_bh30_ch17_0(19); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w65_8 <= DSP_bh30_ch17_0(18); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w64_9 <= DSP_bh30_ch17_0(17); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w63_8 <= DSP_bh30_ch17_0(16); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w62_7 <= DSP_bh30_ch17_0(15); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w61_8 <= DSP_bh30_ch17_0(14); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w60_8 <= DSP_bh30_ch17_0(13); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w59_7 <= DSP_bh30_ch17_0(12); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w58_8 <= DSP_bh30_ch17_0(11); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w57_8 <= DSP_bh30_ch17_0(10); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w56_7 <= DSP_bh30_ch17_0(9); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w55_8 <= DSP_bh30_ch17_0(8); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w54_8 <= DSP_bh30_ch17_0(7); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w53_7 <= DSP_bh30_ch17_0(6); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w52_8 <= DSP_bh30_ch17_0(5); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w51_8 <= DSP_bh30_ch17_0(4); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w50_7 <= DSP_bh30_ch17_0(3); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w49_7 <= DSP_bh30_ch17_0(2); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w48_7 <= DSP_bh30_ch17_0(1); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w47_6 <= DSP_bh30_ch17_0(0); -- cycle= 0 cp= 2.387e-09
   DSP_bh30_ch18_0 <= std_logic_vector(unsigned("" & XX_m29(41 downto 18) & "") * unsigned("" & YY_m29(21 downto 5) & ""));
   heap_bh30_w63_9 <= DSP_bh30_ch18_0(40); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w62_8 <= DSP_bh30_ch18_0(39); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w61_9 <= DSP_bh30_ch18_0(38); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w60_9 <= DSP_bh30_ch18_0(37); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w59_8 <= DSP_bh30_ch18_0(36); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w58_9 <= DSP_bh30_ch18_0(35); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w57_9 <= DSP_bh30_ch18_0(34); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w56_8 <= DSP_bh30_ch18_0(33); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w55_9 <= DSP_bh30_ch18_0(32); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w54_9 <= DSP_bh30_ch18_0(31); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w53_8 <= DSP_bh30_ch18_0(30); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w52_9 <= DSP_bh30_ch18_0(29); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w51_9 <= DSP_bh30_ch18_0(28); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w50_8 <= DSP_bh30_ch18_0(27); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w49_8 <= DSP_bh30_ch18_0(26); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w48_8 <= DSP_bh30_ch18_0(25); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w47_7 <= DSP_bh30_ch18_0(24); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w46_7 <= DSP_bh30_ch18_0(23); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w45_7 <= DSP_bh30_ch18_0(22); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w44_6 <= DSP_bh30_ch18_0(21); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w43_7 <= DSP_bh30_ch18_0(20); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w42_7 <= DSP_bh30_ch18_0(19); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w41_6 <= DSP_bh30_ch18_0(18); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w40_7 <= DSP_bh30_ch18_0(17); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w39_6 <= DSP_bh30_ch18_0(16); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w38_5 <= DSP_bh30_ch18_0(15); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w37_6 <= DSP_bh30_ch18_0(14); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w36_6 <= DSP_bh30_ch18_0(13); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w35_5 <= DSP_bh30_ch18_0(12); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w34_6 <= DSP_bh30_ch18_0(11); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w33_6 <= DSP_bh30_ch18_0(10); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w32_4 <= DSP_bh30_ch18_0(9); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w31_5 <= DSP_bh30_ch18_0(8); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w30_5 <= DSP_bh30_ch18_0(7); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w29_4 <= DSP_bh30_ch18_0(6); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w28_5 <= DSP_bh30_ch18_0(5); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w27_5 <= DSP_bh30_ch18_0(4); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w26_4 <= DSP_bh30_ch18_0(3); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w25_5 <= DSP_bh30_ch18_0(2); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w24_5 <= DSP_bh30_ch18_0(1); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w23_4 <= DSP_bh30_ch18_0(0); -- cycle= 0 cp= 2.387e-09
   DSP_bh30_ch19_0 <= std_logic_vector(unsigned("" & XX_m29(17 downto 0) & "000000") * unsigned("" & YY_m29(21 downto 5) & ""));
   heap_bh30_w39_7 <= DSP_bh30_ch19_0(40); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w38_6 <= DSP_bh30_ch19_0(39); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w37_7 <= DSP_bh30_ch19_0(38); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w36_7 <= DSP_bh30_ch19_0(37); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w35_6 <= DSP_bh30_ch19_0(36); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w34_7 <= DSP_bh30_ch19_0(35); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w33_7 <= DSP_bh30_ch19_0(34); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w32_5 <= DSP_bh30_ch19_0(33); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w31_6 <= DSP_bh30_ch19_0(32); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w30_6 <= DSP_bh30_ch19_0(31); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w29_5 <= DSP_bh30_ch19_0(30); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w28_6 <= DSP_bh30_ch19_0(29); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w27_6 <= DSP_bh30_ch19_0(28); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w26_5 <= DSP_bh30_ch19_0(27); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w25_6 <= DSP_bh30_ch19_0(26); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w24_6 <= DSP_bh30_ch19_0(25); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w23_5 <= DSP_bh30_ch19_0(24); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w22_5 <= DSP_bh30_ch19_0(23); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w21_5 <= DSP_bh30_ch19_0(22); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w20_4 <= DSP_bh30_ch19_0(21); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w19_5 <= DSP_bh30_ch19_0(20); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w18_5 <= DSP_bh30_ch19_0(19); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w17_4 <= DSP_bh30_ch19_0(18); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w16_5 <= DSP_bh30_ch19_0(17); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w15_4 <= DSP_bh30_ch19_0(16); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w14_3 <= DSP_bh30_ch19_0(15); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w13_4 <= DSP_bh30_ch19_0(14); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w12_4 <= DSP_bh30_ch19_0(13); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w11_3 <= DSP_bh30_ch19_0(12); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w10_4 <= DSP_bh30_ch19_0(11); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w9_4 <= DSP_bh30_ch19_0(10); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w8_3 <= DSP_bh30_ch19_0(9); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w7_4 <= DSP_bh30_ch19_0(8); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w6_4 <= DSP_bh30_ch19_0(7); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w5_3 <= DSP_bh30_ch19_0(6); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w4_3 <= DSP_bh30_ch19_0(5); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w3_3 <= DSP_bh30_ch19_0(4); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w2_2 <= DSP_bh30_ch19_0(3); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w1_1 <= DSP_bh30_ch19_0(2); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w0_1 <= DSP_bh30_ch19_0(1); -- cycle= 0 cp= 2.387e-09

   -- Adding the constant bits
      -- All the constant bits are zero, nothing to add


   CompressorIn_bh30_0_0 <= heap_bh30_w6_3 & heap_bh30_w6_2 & heap_bh30_w6_1 & heap_bh30_w6_0;
   CompressorIn_bh30_0_1(0) <= heap_bh30_w7_3;
      Compressor_bh30_0: Compressor_14_3
      port map ( R => CompressorOut_bh30_0_0,
                 X0 => CompressorIn_bh30_0_0,
                 X1 => CompressorIn_bh30_0_1);
   heap_bh30_w6_5 <= CompressorOut_bh30_0_0(0); -- cycle= 0 cp= 1.10504e-09
   heap_bh30_w7_5 <= CompressorOut_bh30_0_0(1); -- cycle= 0 cp= 1.10504e-09
   heap_bh30_w8_4 <= CompressorOut_bh30_0_0(2); -- cycle= 0 cp= 1.10504e-09

   CompressorIn_bh30_1_2 <= heap_bh30_w9_3 & heap_bh30_w9_2 & heap_bh30_w9_1 & heap_bh30_w9_0;
   CompressorIn_bh30_1_3(0) <= heap_bh30_w10_3;
      Compressor_bh30_1: Compressor_14_3
      port map ( R => CompressorOut_bh30_1_1,
                 X0 => CompressorIn_bh30_1_2,
                 X1 => CompressorIn_bh30_1_3);
   heap_bh30_w9_5 <= CompressorOut_bh30_1_1(0); -- cycle= 0 cp= 1.10504e-09
   heap_bh30_w10_5 <= CompressorOut_bh30_1_1(1); -- cycle= 0 cp= 1.10504e-09
   heap_bh30_w11_4 <= CompressorOut_bh30_1_1(2); -- cycle= 0 cp= 1.10504e-09

   CompressorIn_bh30_2_4 <= heap_bh30_w12_3 & heap_bh30_w12_2 & heap_bh30_w12_1 & heap_bh30_w12_0;
   CompressorIn_bh30_2_5(0) <= heap_bh30_w13_3;
      Compressor_bh30_2: Compressor_14_3
      port map ( R => CompressorOut_bh30_2_2,
                 X0 => CompressorIn_bh30_2_4,
                 X1 => CompressorIn_bh30_2_5);
   heap_bh30_w12_5 <= CompressorOut_bh30_2_2(0); -- cycle= 0 cp= 1.10504e-09
   heap_bh30_w13_5 <= CompressorOut_bh30_2_2(1); -- cycle= 0 cp= 1.10504e-09
   heap_bh30_w14_4 <= CompressorOut_bh30_2_2(2); -- cycle= 0 cp= 1.10504e-09

   CompressorIn_bh30_3_6 <= heap_bh30_w15_3 & heap_bh30_w15_2 & heap_bh30_w15_1 & heap_bh30_w15_0;
   CompressorIn_bh30_3_7(0) <= heap_bh30_w16_3;
      Compressor_bh30_3: Compressor_14_3
      port map ( R => CompressorOut_bh30_3_3,
                 X0 => CompressorIn_bh30_3_6,
                 X1 => CompressorIn_bh30_3_7);
   heap_bh30_w15_5 <= CompressorOut_bh30_3_3(0); -- cycle= 0 cp= 1.10504e-09
   heap_bh30_w16_6 <= CompressorOut_bh30_3_3(1); -- cycle= 0 cp= 1.10504e-09
   heap_bh30_w17_5 <= CompressorOut_bh30_3_3(2); -- cycle= 0 cp= 1.10504e-09

   CompressorIn_bh30_4_8 <= heap_bh30_w18_3 & heap_bh30_w18_2 & heap_bh30_w18_1 & heap_bh30_w18_0;
   CompressorIn_bh30_4_9(0) <= heap_bh30_w19_3;
      Compressor_bh30_4: Compressor_14_3
      port map ( R => CompressorOut_bh30_4_4,
                 X0 => CompressorIn_bh30_4_8,
                 X1 => CompressorIn_bh30_4_9);
   heap_bh30_w18_6 <= CompressorOut_bh30_4_4(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w19_6 <= CompressorOut_bh30_4_4(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w20_5 <= CompressorOut_bh30_4_4(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_5_10 <= heap_bh30_w21_3 & heap_bh30_w21_2 & heap_bh30_w21_1 & heap_bh30_w21_0;
   CompressorIn_bh30_5_11(0) <= heap_bh30_w22_3;
      Compressor_bh30_5: Compressor_14_3
      port map ( R => CompressorOut_bh30_5_5,
                 X0 => CompressorIn_bh30_5_10,
                 X1 => CompressorIn_bh30_5_11);
   heap_bh30_w21_6 <= CompressorOut_bh30_5_5(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w22_6 <= CompressorOut_bh30_5_5(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w23_6 <= CompressorOut_bh30_5_5(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_6_12 <= heap_bh30_w24_3 & heap_bh30_w24_2 & heap_bh30_w24_1 & heap_bh30_w24_0;
   CompressorIn_bh30_6_13(0) <= heap_bh30_w25_3;
      Compressor_bh30_6: Compressor_14_3
      port map ( R => CompressorOut_bh30_6_6,
                 X0 => CompressorIn_bh30_6_12,
                 X1 => CompressorIn_bh30_6_13);
   heap_bh30_w24_7 <= CompressorOut_bh30_6_6(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w25_7 <= CompressorOut_bh30_6_6(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w26_6 <= CompressorOut_bh30_6_6(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_7_14 <= heap_bh30_w27_3 & heap_bh30_w27_2 & heap_bh30_w27_1 & heap_bh30_w27_0;
   CompressorIn_bh30_7_15(0) <= heap_bh30_w28_3;
      Compressor_bh30_7: Compressor_14_3
      port map ( R => CompressorOut_bh30_7_7,
                 X0 => CompressorIn_bh30_7_14,
                 X1 => CompressorIn_bh30_7_15);
   heap_bh30_w27_7 <= CompressorOut_bh30_7_7(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w28_7 <= CompressorOut_bh30_7_7(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w29_6 <= CompressorOut_bh30_7_7(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_8_16 <= heap_bh30_w30_3 & heap_bh30_w30_2 & heap_bh30_w30_1 & heap_bh30_w30_0;
   CompressorIn_bh30_8_17(0) <= heap_bh30_w31_3;
      Compressor_bh30_8: Compressor_14_3
      port map ( R => CompressorOut_bh30_8_8,
                 X0 => CompressorIn_bh30_8_16,
                 X1 => CompressorIn_bh30_8_17);
   heap_bh30_w30_7 <= CompressorOut_bh30_8_8(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w31_7 <= CompressorOut_bh30_8_8(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w32_6 <= CompressorOut_bh30_8_8(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_9_18 <= heap_bh30_w33_3 & heap_bh30_w33_2 & heap_bh30_w33_1 & heap_bh30_w33_0;
   CompressorIn_bh30_9_19(0) <= heap_bh30_w34_3;
      Compressor_bh30_9: Compressor_14_3
      port map ( R => CompressorOut_bh30_9_9,
                 X0 => CompressorIn_bh30_9_18,
                 X1 => CompressorIn_bh30_9_19);
   heap_bh30_w33_8 <= CompressorOut_bh30_9_9(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w34_8 <= CompressorOut_bh30_9_9(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w35_7 <= CompressorOut_bh30_9_9(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_10_20 <= heap_bh30_w36_3 & heap_bh30_w36_2 & heap_bh30_w36_1 & heap_bh30_w36_0;
   CompressorIn_bh30_10_21(0) <= heap_bh30_w37_3;
      Compressor_bh30_10: Compressor_14_3
      port map ( R => CompressorOut_bh30_10_10,
                 X0 => CompressorIn_bh30_10_20,
                 X1 => CompressorIn_bh30_10_21);
   heap_bh30_w36_8 <= CompressorOut_bh30_10_10(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w37_8 <= CompressorOut_bh30_10_10(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w38_7 <= CompressorOut_bh30_10_10(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_11_22 <= heap_bh30_w39_3 & heap_bh30_w39_2 & heap_bh30_w39_1 & heap_bh30_w39_0;
   CompressorIn_bh30_11_23(0) <= heap_bh30_w40_3;
      Compressor_bh30_11: Compressor_14_3
      port map ( R => CompressorOut_bh30_11_11,
                 X0 => CompressorIn_bh30_11_22,
                 X1 => CompressorIn_bh30_11_23);
   heap_bh30_w39_8 <= CompressorOut_bh30_11_11(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w40_8 <= CompressorOut_bh30_11_11(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w41_7 <= CompressorOut_bh30_11_11(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_12_24 <= heap_bh30_w42_3 & heap_bh30_w42_2 & heap_bh30_w42_1 & heap_bh30_w42_0;
   CompressorIn_bh30_12_25(0) <= heap_bh30_w43_3;
      Compressor_bh30_12: Compressor_14_3
      port map ( R => CompressorOut_bh30_12_12,
                 X0 => CompressorIn_bh30_12_24,
                 X1 => CompressorIn_bh30_12_25);
   heap_bh30_w42_8 <= CompressorOut_bh30_12_12(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w43_8 <= CompressorOut_bh30_12_12(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w44_7 <= CompressorOut_bh30_12_12(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_13_26 <= heap_bh30_w45_3 & heap_bh30_w45_2 & heap_bh30_w45_1 & heap_bh30_w45_0;
   CompressorIn_bh30_13_27(0) <= heap_bh30_w46_3;
      Compressor_bh30_13: Compressor_14_3
      port map ( R => CompressorOut_bh30_13_13,
                 X0 => CompressorIn_bh30_13_26,
                 X1 => CompressorIn_bh30_13_27);
   heap_bh30_w45_8 <= CompressorOut_bh30_13_13(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w46_8 <= CompressorOut_bh30_13_13(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w47_8 <= CompressorOut_bh30_13_13(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_14_28 <= heap_bh30_w48_3 & heap_bh30_w48_2 & heap_bh30_w48_1 & heap_bh30_w48_0;
   CompressorIn_bh30_14_29(0) <= heap_bh30_w49_3;
      Compressor_bh30_14: Compressor_14_3
      port map ( R => CompressorOut_bh30_14_14,
                 X0 => CompressorIn_bh30_14_28,
                 X1 => CompressorIn_bh30_14_29);
   heap_bh30_w48_9 <= CompressorOut_bh30_14_14(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w49_9 <= CompressorOut_bh30_14_14(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w50_9 <= CompressorOut_bh30_14_14(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_15_30 <= heap_bh30_w51_3 & heap_bh30_w51_2 & heap_bh30_w51_1 & heap_bh30_w51_0;
   CompressorIn_bh30_15_31(0) <= heap_bh30_w52_3;
      Compressor_bh30_15: Compressor_14_3
      port map ( R => CompressorOut_bh30_15_15,
                 X0 => CompressorIn_bh30_15_30,
                 X1 => CompressorIn_bh30_15_31);
   heap_bh30_w51_10 <= CompressorOut_bh30_15_15(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w52_10 <= CompressorOut_bh30_15_15(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w53_9 <= CompressorOut_bh30_15_15(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_16_32 <= heap_bh30_w54_3 & heap_bh30_w54_2 & heap_bh30_w54_1 & heap_bh30_w54_0;
   CompressorIn_bh30_16_33(0) <= heap_bh30_w55_3;
      Compressor_bh30_16: Compressor_14_3
      port map ( R => CompressorOut_bh30_16_16,
                 X0 => CompressorIn_bh30_16_32,
                 X1 => CompressorIn_bh30_16_33);
   heap_bh30_w54_10 <= CompressorOut_bh30_16_16(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w55_10 <= CompressorOut_bh30_16_16(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w56_9 <= CompressorOut_bh30_16_16(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_17_34 <= heap_bh30_w57_3 & heap_bh30_w57_2 & heap_bh30_w57_1 & heap_bh30_w57_0;
   CompressorIn_bh30_17_35(0) <= heap_bh30_w58_3;
      Compressor_bh30_17: Compressor_14_3
      port map ( R => CompressorOut_bh30_17_17,
                 X0 => CompressorIn_bh30_17_34,
                 X1 => CompressorIn_bh30_17_35);
   heap_bh30_w57_10 <= CompressorOut_bh30_17_17(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w58_10 <= CompressorOut_bh30_17_17(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w59_9 <= CompressorOut_bh30_17_17(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_18_36 <= heap_bh30_w60_3 & heap_bh30_w60_2 & heap_bh30_w60_1 & heap_bh30_w60_0;
   CompressorIn_bh30_18_37(0) <= heap_bh30_w61_3;
      Compressor_bh30_18: Compressor_14_3
      port map ( R => CompressorOut_bh30_18_18,
                 X0 => CompressorIn_bh30_18_36,
                 X1 => CompressorIn_bh30_18_37);
   heap_bh30_w60_10 <= CompressorOut_bh30_18_18(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w61_10 <= CompressorOut_bh30_18_18(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w62_9 <= CompressorOut_bh30_18_18(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_19_38 <= heap_bh30_w63_3 & heap_bh30_w63_2 & heap_bh30_w63_1 & heap_bh30_w63_0;
   CompressorIn_bh30_19_39(0) <= heap_bh30_w64_3;
      Compressor_bh30_19: Compressor_14_3
      port map ( R => CompressorOut_bh30_19_19,
                 X0 => CompressorIn_bh30_19_38,
                 X1 => CompressorIn_bh30_19_39);
   heap_bh30_w63_10 <= CompressorOut_bh30_19_19(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w64_10 <= CompressorOut_bh30_19_19(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w65_9 <= CompressorOut_bh30_19_19(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_20_40 <= heap_bh30_w66_3 & heap_bh30_w66_2 & heap_bh30_w66_1 & heap_bh30_w66_0;
   CompressorIn_bh30_20_41(0) <= heap_bh30_w67_3;
      Compressor_bh30_20: Compressor_14_3
      port map ( R => CompressorOut_bh30_20_20,
                 X0 => CompressorIn_bh30_20_40,
                 X1 => CompressorIn_bh30_20_41);
   heap_bh30_w66_10 <= CompressorOut_bh30_20_20(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w67_11 <= CompressorOut_bh30_20_20(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w68_10 <= CompressorOut_bh30_20_20(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_21_42 <= heap_bh30_w69_3 & heap_bh30_w69_2 & heap_bh30_w69_1 & heap_bh30_w69_0;
   CompressorIn_bh30_21_43(0) <= heap_bh30_w70_3;
      Compressor_bh30_21: Compressor_14_3
      port map ( R => CompressorOut_bh30_21_21,
                 X0 => CompressorIn_bh30_21_42,
                 X1 => CompressorIn_bh30_21_43);
   heap_bh30_w69_11 <= CompressorOut_bh30_21_21(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w70_11 <= CompressorOut_bh30_21_21(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w71_11 <= CompressorOut_bh30_21_21(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_22_44 <= heap_bh30_w72_3 & heap_bh30_w72_2 & heap_bh30_w72_1 & heap_bh30_w72_0;
   CompressorIn_bh30_22_45(0) <= heap_bh30_w73_3;
      Compressor_bh30_22: Compressor_14_3
      port map ( R => CompressorOut_bh30_22_22,
                 X0 => CompressorIn_bh30_22_44,
                 X1 => CompressorIn_bh30_22_45);
   heap_bh30_w72_12 <= CompressorOut_bh30_22_22(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w73_12 <= CompressorOut_bh30_22_22(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w74_11 <= CompressorOut_bh30_22_22(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_23_46 <= heap_bh30_w75_3 & heap_bh30_w75_2 & heap_bh30_w75_1 & heap_bh30_w75_0;
   CompressorIn_bh30_23_47(0) <= heap_bh30_w76_3;
      Compressor_bh30_23: Compressor_14_3
      port map ( R => CompressorOut_bh30_23_23,
                 X0 => CompressorIn_bh30_23_46,
                 X1 => CompressorIn_bh30_23_47);
   heap_bh30_w75_12 <= CompressorOut_bh30_23_23(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w76_12 <= CompressorOut_bh30_23_23(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w77_11 <= CompressorOut_bh30_23_23(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_24_48 <= heap_bh30_w78_3 & heap_bh30_w78_2 & heap_bh30_w78_1 & heap_bh30_w78_0;
   CompressorIn_bh30_24_49(0) <= heap_bh30_w79_3;
      Compressor_bh30_24: Compressor_14_3
      port map ( R => CompressorOut_bh30_24_24,
                 X0 => CompressorIn_bh30_24_48,
                 X1 => CompressorIn_bh30_24_49);
   heap_bh30_w78_12 <= CompressorOut_bh30_24_24(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w79_12 <= CompressorOut_bh30_24_24(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w80_11 <= CompressorOut_bh30_24_24(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_25_50 <= heap_bh30_w81_3 & heap_bh30_w81_2 & heap_bh30_w81_1 & heap_bh30_w81_0;
   CompressorIn_bh30_25_51(0) <= heap_bh30_w82_3;
      Compressor_bh30_25: Compressor_14_3
      port map ( R => CompressorOut_bh30_25_25,
                 X0 => CompressorIn_bh30_25_50,
                 X1 => CompressorIn_bh30_25_51);
   heap_bh30_w81_12 <= CompressorOut_bh30_25_25(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w82_12 <= CompressorOut_bh30_25_25(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w83_11 <= CompressorOut_bh30_25_25(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_26_52 <= heap_bh30_w84_3 & heap_bh30_w84_2 & heap_bh30_w84_1 & heap_bh30_w84_0;
   CompressorIn_bh30_26_53(0) <= heap_bh30_w85_3;
      Compressor_bh30_26: Compressor_14_3
      port map ( R => CompressorOut_bh30_26_26,
                 X0 => CompressorIn_bh30_26_52,
                 X1 => CompressorIn_bh30_26_53);
   heap_bh30_w84_12 <= CompressorOut_bh30_26_26(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w85_12 <= CompressorOut_bh30_26_26(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w86_11 <= CompressorOut_bh30_26_26(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_27_54 <= heap_bh30_w87_3 & heap_bh30_w87_2 & heap_bh30_w87_1 & heap_bh30_w87_0;
   CompressorIn_bh30_27_55(0) <= heap_bh30_w88_3;
      Compressor_bh30_27: Compressor_14_3
      port map ( R => CompressorOut_bh30_27_27,
                 X0 => CompressorIn_bh30_27_54,
                 X1 => CompressorIn_bh30_27_55);
   heap_bh30_w87_12 <= CompressorOut_bh30_27_27(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w88_12 <= CompressorOut_bh30_27_27(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w89_11 <= CompressorOut_bh30_27_27(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_28_56 <= heap_bh30_w3_2 & heap_bh30_w3_1 & heap_bh30_w3_0;
   CompressorIn_bh30_28_57 <= heap_bh30_w4_2 & heap_bh30_w4_1;
      Compressor_bh30_28: Compressor_23_3
      port map ( R => CompressorOut_bh30_28_28,
                 X0 => CompressorIn_bh30_28_56,
                 X1 => CompressorIn_bh30_28_57);
   heap_bh30_w3_4 <= CompressorOut_bh30_28_28(0); -- cycle= 0 cp= 1.10504e-09
   heap_bh30_w4_4 <= CompressorOut_bh30_28_28(1); -- cycle= 0 cp= 1.10504e-09
   heap_bh30_w5_4 <= CompressorOut_bh30_28_28(2); -- cycle= 0 cp= 1.10504e-09

   CompressorIn_bh30_29_58 <= heap_bh30_w7_2 & heap_bh30_w7_1 & heap_bh30_w7_0;
   CompressorIn_bh30_29_59 <= heap_bh30_w8_2 & heap_bh30_w8_1;
      Compressor_bh30_29: Compressor_23_3
      port map ( R => CompressorOut_bh30_29_29,
                 X0 => CompressorIn_bh30_29_58,
                 X1 => CompressorIn_bh30_29_59);
   heap_bh30_w7_6 <= CompressorOut_bh30_29_29(0); -- cycle= 0 cp= 1.10504e-09
   heap_bh30_w8_5 <= CompressorOut_bh30_29_29(1); -- cycle= 0 cp= 1.10504e-09
   heap_bh30_w9_6 <= CompressorOut_bh30_29_29(2); -- cycle= 0 cp= 1.10504e-09

   CompressorIn_bh30_30_60 <= heap_bh30_w10_2 & heap_bh30_w10_1 & heap_bh30_w10_0;
   CompressorIn_bh30_30_61 <= heap_bh30_w11_2 & heap_bh30_w11_1;
      Compressor_bh30_30: Compressor_23_3
      port map ( R => CompressorOut_bh30_30_30,
                 X0 => CompressorIn_bh30_30_60,
                 X1 => CompressorIn_bh30_30_61);
   heap_bh30_w10_6 <= CompressorOut_bh30_30_30(0); -- cycle= 0 cp= 1.10504e-09
   heap_bh30_w11_5 <= CompressorOut_bh30_30_30(1); -- cycle= 0 cp= 1.10504e-09
   heap_bh30_w12_6 <= CompressorOut_bh30_30_30(2); -- cycle= 0 cp= 1.10504e-09

   CompressorIn_bh30_31_62 <= heap_bh30_w13_2 & heap_bh30_w13_1 & heap_bh30_w13_0;
   CompressorIn_bh30_31_63 <= heap_bh30_w14_2 & heap_bh30_w14_1;
      Compressor_bh30_31: Compressor_23_3
      port map ( R => CompressorOut_bh30_31_31,
                 X0 => CompressorIn_bh30_31_62,
                 X1 => CompressorIn_bh30_31_63);
   heap_bh30_w13_6 <= CompressorOut_bh30_31_31(0); -- cycle= 0 cp= 1.10504e-09
   heap_bh30_w14_5 <= CompressorOut_bh30_31_31(1); -- cycle= 0 cp= 1.10504e-09
   heap_bh30_w15_6 <= CompressorOut_bh30_31_31(2); -- cycle= 0 cp= 1.10504e-09

   CompressorIn_bh30_32_64 <= heap_bh30_w16_2 & heap_bh30_w16_1 & heap_bh30_w16_0;
   CompressorIn_bh30_32_65 <= heap_bh30_w17_2 & heap_bh30_w17_1;
      Compressor_bh30_32: Compressor_23_3
      port map ( R => CompressorOut_bh30_32_32,
                 X0 => CompressorIn_bh30_32_64,
                 X1 => CompressorIn_bh30_32_65);
   heap_bh30_w16_7 <= CompressorOut_bh30_32_32(0); -- cycle= 0 cp= 1.10504e-09
   heap_bh30_w17_6 <= CompressorOut_bh30_32_32(1); -- cycle= 0 cp= 1.10504e-09
   heap_bh30_w18_7 <= CompressorOut_bh30_32_32(2); -- cycle= 0 cp= 1.10504e-09

   CompressorIn_bh30_33_66 <= heap_bh30_w19_2 & heap_bh30_w19_1 & heap_bh30_w19_0;
   CompressorIn_bh30_33_67 <= heap_bh30_w20_2 & heap_bh30_w20_1;
      Compressor_bh30_33: Compressor_23_3
      port map ( R => CompressorOut_bh30_33_33,
                 X0 => CompressorIn_bh30_33_66,
                 X1 => CompressorIn_bh30_33_67);
   heap_bh30_w19_7 <= CompressorOut_bh30_33_33(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w20_6 <= CompressorOut_bh30_33_33(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w21_7 <= CompressorOut_bh30_33_33(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_34_68 <= heap_bh30_w22_2 & heap_bh30_w22_1 & heap_bh30_w22_0;
   CompressorIn_bh30_34_69 <= heap_bh30_w23_2 & heap_bh30_w23_1;
      Compressor_bh30_34: Compressor_23_3
      port map ( R => CompressorOut_bh30_34_34,
                 X0 => CompressorIn_bh30_34_68,
                 X1 => CompressorIn_bh30_34_69);
   heap_bh30_w22_7 <= CompressorOut_bh30_34_34(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w23_7 <= CompressorOut_bh30_34_34(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w24_8 <= CompressorOut_bh30_34_34(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_35_70 <= heap_bh30_w25_2 & heap_bh30_w25_1 & heap_bh30_w25_0;
   CompressorIn_bh30_35_71 <= heap_bh30_w26_2 & heap_bh30_w26_1;
      Compressor_bh30_35: Compressor_23_3
      port map ( R => CompressorOut_bh30_35_35,
                 X0 => CompressorIn_bh30_35_70,
                 X1 => CompressorIn_bh30_35_71);
   heap_bh30_w25_8 <= CompressorOut_bh30_35_35(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w26_7 <= CompressorOut_bh30_35_35(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w27_8 <= CompressorOut_bh30_35_35(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_36_72 <= heap_bh30_w28_2 & heap_bh30_w28_1 & heap_bh30_w28_0;
   CompressorIn_bh30_36_73 <= heap_bh30_w29_2 & heap_bh30_w29_1;
      Compressor_bh30_36: Compressor_23_3
      port map ( R => CompressorOut_bh30_36_36,
                 X0 => CompressorIn_bh30_36_72,
                 X1 => CompressorIn_bh30_36_73);
   heap_bh30_w28_8 <= CompressorOut_bh30_36_36(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w29_7 <= CompressorOut_bh30_36_36(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w30_8 <= CompressorOut_bh30_36_36(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_37_74 <= heap_bh30_w31_2 & heap_bh30_w31_1 & heap_bh30_w31_0;
   CompressorIn_bh30_37_75 <= heap_bh30_w32_2 & heap_bh30_w32_1;
      Compressor_bh30_37: Compressor_23_3
      port map ( R => CompressorOut_bh30_37_37,
                 X0 => CompressorIn_bh30_37_74,
                 X1 => CompressorIn_bh30_37_75);
   heap_bh30_w31_8 <= CompressorOut_bh30_37_37(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w32_7 <= CompressorOut_bh30_37_37(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w33_9 <= CompressorOut_bh30_37_37(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_38_76 <= heap_bh30_w34_2 & heap_bh30_w34_1 & heap_bh30_w34_0;
   CompressorIn_bh30_38_77 <= heap_bh30_w35_2 & heap_bh30_w35_1;
      Compressor_bh30_38: Compressor_23_3
      port map ( R => CompressorOut_bh30_38_38,
                 X0 => CompressorIn_bh30_38_76,
                 X1 => CompressorIn_bh30_38_77);
   heap_bh30_w34_9 <= CompressorOut_bh30_38_38(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w35_8 <= CompressorOut_bh30_38_38(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w36_9 <= CompressorOut_bh30_38_38(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_39_78 <= heap_bh30_w37_2 & heap_bh30_w37_1 & heap_bh30_w37_0;
   CompressorIn_bh30_39_79 <= heap_bh30_w38_2 & heap_bh30_w38_1;
      Compressor_bh30_39: Compressor_23_3
      port map ( R => CompressorOut_bh30_39_39,
                 X0 => CompressorIn_bh30_39_78,
                 X1 => CompressorIn_bh30_39_79);
   heap_bh30_w37_9 <= CompressorOut_bh30_39_39(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w38_8 <= CompressorOut_bh30_39_39(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w39_9 <= CompressorOut_bh30_39_39(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_40_80 <= heap_bh30_w40_2 & heap_bh30_w40_1 & heap_bh30_w40_0;
   CompressorIn_bh30_40_81 <= heap_bh30_w41_2 & heap_bh30_w41_1;
      Compressor_bh30_40: Compressor_23_3
      port map ( R => CompressorOut_bh30_40_40,
                 X0 => CompressorIn_bh30_40_80,
                 X1 => CompressorIn_bh30_40_81);
   heap_bh30_w40_9 <= CompressorOut_bh30_40_40(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w41_8 <= CompressorOut_bh30_40_40(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w42_9 <= CompressorOut_bh30_40_40(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_41_82 <= heap_bh30_w43_2 & heap_bh30_w43_1 & heap_bh30_w43_0;
   CompressorIn_bh30_41_83 <= heap_bh30_w44_2 & heap_bh30_w44_1;
      Compressor_bh30_41: Compressor_23_3
      port map ( R => CompressorOut_bh30_41_41,
                 X0 => CompressorIn_bh30_41_82,
                 X1 => CompressorIn_bh30_41_83);
   heap_bh30_w43_9 <= CompressorOut_bh30_41_41(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w44_8 <= CompressorOut_bh30_41_41(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w45_9 <= CompressorOut_bh30_41_41(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_42_84 <= heap_bh30_w46_2 & heap_bh30_w46_1 & heap_bh30_w46_0;
   CompressorIn_bh30_42_85 <= heap_bh30_w47_2 & heap_bh30_w47_1;
      Compressor_bh30_42: Compressor_23_3
      port map ( R => CompressorOut_bh30_42_42,
                 X0 => CompressorIn_bh30_42_84,
                 X1 => CompressorIn_bh30_42_85);
   heap_bh30_w46_9 <= CompressorOut_bh30_42_42(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w47_9 <= CompressorOut_bh30_42_42(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w48_10 <= CompressorOut_bh30_42_42(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_43_86 <= heap_bh30_w49_2 & heap_bh30_w49_1 & heap_bh30_w49_0;
   CompressorIn_bh30_43_87 <= heap_bh30_w50_2 & heap_bh30_w50_1;
      Compressor_bh30_43: Compressor_23_3
      port map ( R => CompressorOut_bh30_43_43,
                 X0 => CompressorIn_bh30_43_86,
                 X1 => CompressorIn_bh30_43_87);
   heap_bh30_w49_10 <= CompressorOut_bh30_43_43(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w50_10 <= CompressorOut_bh30_43_43(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w51_11 <= CompressorOut_bh30_43_43(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_44_88 <= heap_bh30_w52_2 & heap_bh30_w52_1 & heap_bh30_w52_0;
   CompressorIn_bh30_44_89 <= heap_bh30_w53_2 & heap_bh30_w53_1;
      Compressor_bh30_44: Compressor_23_3
      port map ( R => CompressorOut_bh30_44_44,
                 X0 => CompressorIn_bh30_44_88,
                 X1 => CompressorIn_bh30_44_89);
   heap_bh30_w52_11 <= CompressorOut_bh30_44_44(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w53_10 <= CompressorOut_bh30_44_44(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w54_11 <= CompressorOut_bh30_44_44(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_45_90 <= heap_bh30_w55_2 & heap_bh30_w55_1 & heap_bh30_w55_0;
   CompressorIn_bh30_45_91 <= heap_bh30_w56_2 & heap_bh30_w56_1;
      Compressor_bh30_45: Compressor_23_3
      port map ( R => CompressorOut_bh30_45_45,
                 X0 => CompressorIn_bh30_45_90,
                 X1 => CompressorIn_bh30_45_91);
   heap_bh30_w55_11 <= CompressorOut_bh30_45_45(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w56_10 <= CompressorOut_bh30_45_45(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w57_11 <= CompressorOut_bh30_45_45(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_46_92 <= heap_bh30_w58_2 & heap_bh30_w58_1 & heap_bh30_w58_0;
   CompressorIn_bh30_46_93 <= heap_bh30_w59_2 & heap_bh30_w59_1;
      Compressor_bh30_46: Compressor_23_3
      port map ( R => CompressorOut_bh30_46_46,
                 X0 => CompressorIn_bh30_46_92,
                 X1 => CompressorIn_bh30_46_93);
   heap_bh30_w58_11 <= CompressorOut_bh30_46_46(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w59_10 <= CompressorOut_bh30_46_46(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w60_11 <= CompressorOut_bh30_46_46(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_47_94 <= heap_bh30_w61_2 & heap_bh30_w61_1 & heap_bh30_w61_0;
   CompressorIn_bh30_47_95 <= heap_bh30_w62_2 & heap_bh30_w62_1;
      Compressor_bh30_47: Compressor_23_3
      port map ( R => CompressorOut_bh30_47_47,
                 X0 => CompressorIn_bh30_47_94,
                 X1 => CompressorIn_bh30_47_95);
   heap_bh30_w61_11 <= CompressorOut_bh30_47_47(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w62_10 <= CompressorOut_bh30_47_47(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w63_11 <= CompressorOut_bh30_47_47(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_48_96 <= heap_bh30_w64_2 & heap_bh30_w64_1 & heap_bh30_w64_0;
   CompressorIn_bh30_48_97 <= heap_bh30_w65_2 & heap_bh30_w65_1;
      Compressor_bh30_48: Compressor_23_3
      port map ( R => CompressorOut_bh30_48_48,
                 X0 => CompressorIn_bh30_48_96,
                 X1 => CompressorIn_bh30_48_97);
   heap_bh30_w64_11 <= CompressorOut_bh30_48_48(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w65_10 <= CompressorOut_bh30_48_48(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w66_11 <= CompressorOut_bh30_48_48(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_49_98 <= heap_bh30_w67_2 & heap_bh30_w67_1 & heap_bh30_w67_0;
   CompressorIn_bh30_49_99 <= heap_bh30_w68_2 & heap_bh30_w68_1;
      Compressor_bh30_49: Compressor_23_3
      port map ( R => CompressorOut_bh30_49_49,
                 X0 => CompressorIn_bh30_49_98,
                 X1 => CompressorIn_bh30_49_99);
   heap_bh30_w67_12 <= CompressorOut_bh30_49_49(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w68_11 <= CompressorOut_bh30_49_49(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w69_12 <= CompressorOut_bh30_49_49(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_50_100 <= heap_bh30_w70_2 & heap_bh30_w70_1 & heap_bh30_w70_0;
   CompressorIn_bh30_50_101 <= heap_bh30_w71_2 & heap_bh30_w71_1;
      Compressor_bh30_50: Compressor_23_3
      port map ( R => CompressorOut_bh30_50_50,
                 X0 => CompressorIn_bh30_50_100,
                 X1 => CompressorIn_bh30_50_101);
   heap_bh30_w70_12 <= CompressorOut_bh30_50_50(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w71_12 <= CompressorOut_bh30_50_50(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w72_13 <= CompressorOut_bh30_50_50(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_51_102 <= heap_bh30_w73_2 & heap_bh30_w73_1 & heap_bh30_w73_0;
   CompressorIn_bh30_51_103 <= heap_bh30_w74_2 & heap_bh30_w74_1;
      Compressor_bh30_51: Compressor_23_3
      port map ( R => CompressorOut_bh30_51_51,
                 X0 => CompressorIn_bh30_51_102,
                 X1 => CompressorIn_bh30_51_103);
   heap_bh30_w73_13 <= CompressorOut_bh30_51_51(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w74_12 <= CompressorOut_bh30_51_51(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w75_13 <= CompressorOut_bh30_51_51(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_52_104 <= heap_bh30_w76_2 & heap_bh30_w76_1 & heap_bh30_w76_0;
   CompressorIn_bh30_52_105 <= heap_bh30_w77_2 & heap_bh30_w77_1;
      Compressor_bh30_52: Compressor_23_3
      port map ( R => CompressorOut_bh30_52_52,
                 X0 => CompressorIn_bh30_52_104,
                 X1 => CompressorIn_bh30_52_105);
   heap_bh30_w76_13 <= CompressorOut_bh30_52_52(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w77_12 <= CompressorOut_bh30_52_52(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w78_13 <= CompressorOut_bh30_52_52(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_53_106 <= heap_bh30_w79_2 & heap_bh30_w79_1 & heap_bh30_w79_0;
   CompressorIn_bh30_53_107 <= heap_bh30_w80_2 & heap_bh30_w80_1;
      Compressor_bh30_53: Compressor_23_3
      port map ( R => CompressorOut_bh30_53_53,
                 X0 => CompressorIn_bh30_53_106,
                 X1 => CompressorIn_bh30_53_107);
   heap_bh30_w79_13 <= CompressorOut_bh30_53_53(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w80_12 <= CompressorOut_bh30_53_53(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w81_13 <= CompressorOut_bh30_53_53(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_54_108 <= heap_bh30_w82_2 & heap_bh30_w82_1 & heap_bh30_w82_0;
   CompressorIn_bh30_54_109 <= heap_bh30_w83_2 & heap_bh30_w83_1;
      Compressor_bh30_54: Compressor_23_3
      port map ( R => CompressorOut_bh30_54_54,
                 X0 => CompressorIn_bh30_54_108,
                 X1 => CompressorIn_bh30_54_109);
   heap_bh30_w82_13 <= CompressorOut_bh30_54_54(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w83_12 <= CompressorOut_bh30_54_54(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w84_13 <= CompressorOut_bh30_54_54(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_55_110 <= heap_bh30_w85_2 & heap_bh30_w85_1 & heap_bh30_w85_0;
   CompressorIn_bh30_55_111 <= heap_bh30_w86_2 & heap_bh30_w86_1;
      Compressor_bh30_55: Compressor_23_3
      port map ( R => CompressorOut_bh30_55_55,
                 X0 => CompressorIn_bh30_55_110,
                 X1 => CompressorIn_bh30_55_111);
   heap_bh30_w85_13 <= CompressorOut_bh30_55_55(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w86_12 <= CompressorOut_bh30_55_55(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w87_13 <= CompressorOut_bh30_55_55(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_56_112 <= heap_bh30_w88_2 & heap_bh30_w88_1 & heap_bh30_w88_0;
   CompressorIn_bh30_56_113 <= heap_bh30_w89_2 & heap_bh30_w89_1;
      Compressor_bh30_56: Compressor_23_3
      port map ( R => CompressorOut_bh30_56_56,
                 X0 => CompressorIn_bh30_56_112,
                 X1 => CompressorIn_bh30_56_113);
   heap_bh30_w88_13 <= CompressorOut_bh30_56_56(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w89_12 <= CompressorOut_bh30_56_56(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w90_11 <= CompressorOut_bh30_56_56(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_57_114 <= heap_bh30_w90_2 & heap_bh30_w90_1 & heap_bh30_w90_0;
   CompressorIn_bh30_57_115 <= heap_bh30_w91_2 & heap_bh30_w91_1;
      Compressor_bh30_57: Compressor_23_3
      port map ( R => CompressorOut_bh30_57_57,
                 X0 => CompressorIn_bh30_57_114,
                 X1 => CompressorIn_bh30_57_115);
   heap_bh30_w90_12 <= CompressorOut_bh30_57_57(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w91_11 <= CompressorOut_bh30_57_57(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w92_9 <= CompressorOut_bh30_57_57(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_58_116 <= heap_bh30_w5_2 & heap_bh30_w5_1 & heap_bh30_w5_0;
      Compressor_bh30_58: Compressor_3_2
      port map ( R => CompressorOut_bh30_58_58,
                 X0 => CompressorIn_bh30_58_116);
   heap_bh30_w5_5 <= CompressorOut_bh30_58_58(0); -- cycle= 0 cp= 1.10504e-09
   heap_bh30_w6_6 <= CompressorOut_bh30_58_58(1); -- cycle= 0 cp= 1.10504e-09

   CompressorIn_bh30_59_117 <= heap_bh30_w8_0 & heap_bh30_w8_5 & heap_bh30_w8_4;
   CompressorIn_bh30_59_118 <= heap_bh30_w9_6 & heap_bh30_w9_5;
      Compressor_bh30_59: Compressor_23_3
      port map ( R => CompressorOut_bh30_59_59,
                 X0 => CompressorIn_bh30_59_117,
                 X1 => CompressorIn_bh30_59_118);
   heap_bh30_w8_6 <= CompressorOut_bh30_59_59(0); -- cycle= 0 cp= 1.63576e-09
   heap_bh30_w9_7 <= CompressorOut_bh30_59_59(1); -- cycle= 0 cp= 1.63576e-09
   heap_bh30_w10_7 <= CompressorOut_bh30_59_59(2); -- cycle= 0 cp= 1.63576e-09

   CompressorIn_bh30_60_119 <= heap_bh30_w11_0 & heap_bh30_w11_5 & heap_bh30_w11_4;
   CompressorIn_bh30_60_120 <= heap_bh30_w12_6 & heap_bh30_w12_5;
      Compressor_bh30_60: Compressor_23_3
      port map ( R => CompressorOut_bh30_60_60,
                 X0 => CompressorIn_bh30_60_119,
                 X1 => CompressorIn_bh30_60_120);
   heap_bh30_w11_6 <= CompressorOut_bh30_60_60(0); -- cycle= 0 cp= 1.63576e-09
   heap_bh30_w12_7 <= CompressorOut_bh30_60_60(1); -- cycle= 0 cp= 1.63576e-09
   heap_bh30_w13_7 <= CompressorOut_bh30_60_60(2); -- cycle= 0 cp= 1.63576e-09

   CompressorIn_bh30_61_121 <= heap_bh30_w14_0 & heap_bh30_w14_5 & heap_bh30_w14_4;
   CompressorIn_bh30_61_122 <= heap_bh30_w15_6 & heap_bh30_w15_5;
      Compressor_bh30_61: Compressor_23_3
      port map ( R => CompressorOut_bh30_61_61,
                 X0 => CompressorIn_bh30_61_121,
                 X1 => CompressorIn_bh30_61_122);
   heap_bh30_w14_6 <= CompressorOut_bh30_61_61(0); -- cycle= 0 cp= 1.63576e-09
   heap_bh30_w15_7 <= CompressorOut_bh30_61_61(1); -- cycle= 0 cp= 1.63576e-09
   heap_bh30_w16_8 <= CompressorOut_bh30_61_61(2); -- cycle= 0 cp= 1.63576e-09

   CompressorIn_bh30_62_123 <= heap_bh30_w17_0 & heap_bh30_w17_6 & heap_bh30_w17_5;
   CompressorIn_bh30_62_124 <= heap_bh30_w18_7 & heap_bh30_w18_6;
      Compressor_bh30_62: Compressor_23_3
      port map ( R => CompressorOut_bh30_62_62,
                 X0 => CompressorIn_bh30_62_123,
                 X1 => CompressorIn_bh30_62_124);
   heap_bh30_w17_7 <= CompressorOut_bh30_62_62(0); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w18_8 <= CompressorOut_bh30_62_62(1); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w19_8 <= CompressorOut_bh30_62_62(2); -- cycle= 0 cp= 1.6532e-09

   CompressorIn_bh30_63_125 <= heap_bh30_w20_0 & heap_bh30_w20_6 & heap_bh30_w20_5;
   CompressorIn_bh30_63_126 <= heap_bh30_w21_7 & heap_bh30_w21_6;
      Compressor_bh30_63: Compressor_23_3
      port map ( R => CompressorOut_bh30_63_63,
                 X0 => CompressorIn_bh30_63_125,
                 X1 => CompressorIn_bh30_63_126);
   heap_bh30_w20_7 <= CompressorOut_bh30_63_63(0); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w21_8 <= CompressorOut_bh30_63_63(1); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w22_8 <= CompressorOut_bh30_63_63(2); -- cycle= 0 cp= 1.6532e-09

   CompressorIn_bh30_64_127 <= heap_bh30_w23_0 & heap_bh30_w23_7 & heap_bh30_w23_6;
   CompressorIn_bh30_64_128 <= heap_bh30_w24_8 & heap_bh30_w24_7;
      Compressor_bh30_64: Compressor_23_3
      port map ( R => CompressorOut_bh30_64_64,
                 X0 => CompressorIn_bh30_64_127,
                 X1 => CompressorIn_bh30_64_128);
   heap_bh30_w23_8 <= CompressorOut_bh30_64_64(0); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w24_9 <= CompressorOut_bh30_64_64(1); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w25_9 <= CompressorOut_bh30_64_64(2); -- cycle= 0 cp= 1.6532e-09

   CompressorIn_bh30_65_129 <= heap_bh30_w26_0 & heap_bh30_w26_7 & heap_bh30_w26_6;
   CompressorIn_bh30_65_130 <= heap_bh30_w27_8 & heap_bh30_w27_7;
      Compressor_bh30_65: Compressor_23_3
      port map ( R => CompressorOut_bh30_65_65,
                 X0 => CompressorIn_bh30_65_129,
                 X1 => CompressorIn_bh30_65_130);
   heap_bh30_w26_8 <= CompressorOut_bh30_65_65(0); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w27_9 <= CompressorOut_bh30_65_65(1); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w28_9 <= CompressorOut_bh30_65_65(2); -- cycle= 0 cp= 1.6532e-09

   CompressorIn_bh30_66_131 <= heap_bh30_w29_0 & heap_bh30_w29_7 & heap_bh30_w29_6;
   CompressorIn_bh30_66_132 <= heap_bh30_w30_8 & heap_bh30_w30_7;
      Compressor_bh30_66: Compressor_23_3
      port map ( R => CompressorOut_bh30_66_66,
                 X0 => CompressorIn_bh30_66_131,
                 X1 => CompressorIn_bh30_66_132);
   heap_bh30_w29_8 <= CompressorOut_bh30_66_66(0); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w30_9 <= CompressorOut_bh30_66_66(1); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w31_9 <= CompressorOut_bh30_66_66(2); -- cycle= 0 cp= 1.6532e-09

   CompressorIn_bh30_67_133 <= heap_bh30_w32_0 & heap_bh30_w32_7 & heap_bh30_w32_6;
   CompressorIn_bh30_67_134 <= heap_bh30_w33_9 & heap_bh30_w33_8;
      Compressor_bh30_67: Compressor_23_3
      port map ( R => CompressorOut_bh30_67_67,
                 X0 => CompressorIn_bh30_67_133,
                 X1 => CompressorIn_bh30_67_134);
   heap_bh30_w32_8 <= CompressorOut_bh30_67_67(0); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w33_10 <= CompressorOut_bh30_67_67(1); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w34_10 <= CompressorOut_bh30_67_67(2); -- cycle= 0 cp= 1.6532e-09

   CompressorIn_bh30_68_135 <= heap_bh30_w35_0 & heap_bh30_w35_8 & heap_bh30_w35_7;
   CompressorIn_bh30_68_136 <= heap_bh30_w36_9 & heap_bh30_w36_8;
      Compressor_bh30_68: Compressor_23_3
      port map ( R => CompressorOut_bh30_68_68,
                 X0 => CompressorIn_bh30_68_135,
                 X1 => CompressorIn_bh30_68_136);
   heap_bh30_w35_9 <= CompressorOut_bh30_68_68(0); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w36_10 <= CompressorOut_bh30_68_68(1); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w37_10 <= CompressorOut_bh30_68_68(2); -- cycle= 0 cp= 1.6532e-09

   CompressorIn_bh30_69_137 <= heap_bh30_w38_0 & heap_bh30_w38_8 & heap_bh30_w38_7;
   CompressorIn_bh30_69_138 <= heap_bh30_w39_9 & heap_bh30_w39_8;
      Compressor_bh30_69: Compressor_23_3
      port map ( R => CompressorOut_bh30_69_69,
                 X0 => CompressorIn_bh30_69_137,
                 X1 => CompressorIn_bh30_69_138);
   heap_bh30_w38_9 <= CompressorOut_bh30_69_69(0); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w39_10 <= CompressorOut_bh30_69_69(1); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w40_10 <= CompressorOut_bh30_69_69(2); -- cycle= 0 cp= 1.6532e-09

   CompressorIn_bh30_70_139 <= heap_bh30_w41_0 & heap_bh30_w41_8 & heap_bh30_w41_7;
   CompressorIn_bh30_70_140 <= heap_bh30_w42_9 & heap_bh30_w42_8;
      Compressor_bh30_70: Compressor_23_3
      port map ( R => CompressorOut_bh30_70_70,
                 X0 => CompressorIn_bh30_70_139,
                 X1 => CompressorIn_bh30_70_140);
   heap_bh30_w41_9 <= CompressorOut_bh30_70_70(0); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w42_10 <= CompressorOut_bh30_70_70(1); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w43_10 <= CompressorOut_bh30_70_70(2); -- cycle= 0 cp= 1.6532e-09

   CompressorIn_bh30_71_141 <= heap_bh30_w44_0 & heap_bh30_w44_8 & heap_bh30_w44_7;
   CompressorIn_bh30_71_142 <= heap_bh30_w45_9 & heap_bh30_w45_8;
      Compressor_bh30_71: Compressor_23_3
      port map ( R => CompressorOut_bh30_71_71,
                 X0 => CompressorIn_bh30_71_141,
                 X1 => CompressorIn_bh30_71_142);
   heap_bh30_w44_9 <= CompressorOut_bh30_71_71(0); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w45_10 <= CompressorOut_bh30_71_71(1); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w46_10 <= CompressorOut_bh30_71_71(2); -- cycle= 0 cp= 1.6532e-09

   CompressorIn_bh30_72_143 <= heap_bh30_w47_0 & heap_bh30_w47_9 & heap_bh30_w47_8;
   CompressorIn_bh30_72_144 <= heap_bh30_w48_10 & heap_bh30_w48_9;
      Compressor_bh30_72: Compressor_23_3
      port map ( R => CompressorOut_bh30_72_72,
                 X0 => CompressorIn_bh30_72_143,
                 X1 => CompressorIn_bh30_72_144);
   heap_bh30_w47_10 <= CompressorOut_bh30_72_72(0); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w48_11 <= CompressorOut_bh30_72_72(1); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w49_11 <= CompressorOut_bh30_72_72(2); -- cycle= 0 cp= 1.6532e-09

   CompressorIn_bh30_73_145 <= heap_bh30_w50_0 & heap_bh30_w50_10 & heap_bh30_w50_9;
   CompressorIn_bh30_73_146 <= heap_bh30_w51_11 & heap_bh30_w51_10;
      Compressor_bh30_73: Compressor_23_3
      port map ( R => CompressorOut_bh30_73_73,
                 X0 => CompressorIn_bh30_73_145,
                 X1 => CompressorIn_bh30_73_146);
   heap_bh30_w50_11 <= CompressorOut_bh30_73_73(0); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w51_12 <= CompressorOut_bh30_73_73(1); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w52_12 <= CompressorOut_bh30_73_73(2); -- cycle= 0 cp= 1.6532e-09

   CompressorIn_bh30_74_147 <= heap_bh30_w53_0 & heap_bh30_w53_10 & heap_bh30_w53_9;
   CompressorIn_bh30_74_148 <= heap_bh30_w54_11 & heap_bh30_w54_10;
      Compressor_bh30_74: Compressor_23_3
      port map ( R => CompressorOut_bh30_74_74,
                 X0 => CompressorIn_bh30_74_147,
                 X1 => CompressorIn_bh30_74_148);
   heap_bh30_w53_11 <= CompressorOut_bh30_74_74(0); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w54_12 <= CompressorOut_bh30_74_74(1); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w55_12 <= CompressorOut_bh30_74_74(2); -- cycle= 0 cp= 1.6532e-09

   CompressorIn_bh30_75_149 <= heap_bh30_w56_0 & heap_bh30_w56_10 & heap_bh30_w56_9;
   CompressorIn_bh30_75_150 <= heap_bh30_w57_11 & heap_bh30_w57_10;
      Compressor_bh30_75: Compressor_23_3
      port map ( R => CompressorOut_bh30_75_75,
                 X0 => CompressorIn_bh30_75_149,
                 X1 => CompressorIn_bh30_75_150);
   heap_bh30_w56_11 <= CompressorOut_bh30_75_75(0); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w57_12 <= CompressorOut_bh30_75_75(1); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w58_12 <= CompressorOut_bh30_75_75(2); -- cycle= 0 cp= 1.6532e-09

   CompressorIn_bh30_76_151 <= heap_bh30_w59_0 & heap_bh30_w59_10 & heap_bh30_w59_9;
   CompressorIn_bh30_76_152 <= heap_bh30_w60_11 & heap_bh30_w60_10;
      Compressor_bh30_76: Compressor_23_3
      port map ( R => CompressorOut_bh30_76_76,
                 X0 => CompressorIn_bh30_76_151,
                 X1 => CompressorIn_bh30_76_152);
   heap_bh30_w59_11 <= CompressorOut_bh30_76_76(0); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w60_12 <= CompressorOut_bh30_76_76(1); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w61_12 <= CompressorOut_bh30_76_76(2); -- cycle= 0 cp= 1.6532e-09

   CompressorIn_bh30_77_153 <= heap_bh30_w62_0 & heap_bh30_w62_10 & heap_bh30_w62_9;
   CompressorIn_bh30_77_154 <= heap_bh30_w63_11 & heap_bh30_w63_10;
      Compressor_bh30_77: Compressor_23_3
      port map ( R => CompressorOut_bh30_77_77,
                 X0 => CompressorIn_bh30_77_153,
                 X1 => CompressorIn_bh30_77_154);
   heap_bh30_w62_11 <= CompressorOut_bh30_77_77(0); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w63_12 <= CompressorOut_bh30_77_77(1); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w64_12 <= CompressorOut_bh30_77_77(2); -- cycle= 0 cp= 1.6532e-09

   CompressorIn_bh30_78_155 <= heap_bh30_w65_0 & heap_bh30_w65_10 & heap_bh30_w65_9;
   CompressorIn_bh30_78_156 <= heap_bh30_w66_11 & heap_bh30_w66_10;
      Compressor_bh30_78: Compressor_23_3
      port map ( R => CompressorOut_bh30_78_78,
                 X0 => CompressorIn_bh30_78_155,
                 X1 => CompressorIn_bh30_78_156);
   heap_bh30_w65_11 <= CompressorOut_bh30_78_78(0); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w66_12 <= CompressorOut_bh30_78_78(1); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w67_13 <= CompressorOut_bh30_78_78(2); -- cycle= 0 cp= 1.6532e-09

   CompressorIn_bh30_79_157 <= heap_bh30_w68_0 & heap_bh30_w68_11 & heap_bh30_w68_10;
   CompressorIn_bh30_79_158 <= heap_bh30_w69_12 & heap_bh30_w69_11;
      Compressor_bh30_79: Compressor_23_3
      port map ( R => CompressorOut_bh30_79_79,
                 X0 => CompressorIn_bh30_79_157,
                 X1 => CompressorIn_bh30_79_158);
   heap_bh30_w68_12 <= CompressorOut_bh30_79_79(0); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w69_13 <= CompressorOut_bh30_79_79(1); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w70_13 <= CompressorOut_bh30_79_79(2); -- cycle= 0 cp= 1.6532e-09

   CompressorIn_bh30_80_159 <= heap_bh30_w71_0 & heap_bh30_w71_12 & heap_bh30_w71_11;
   CompressorIn_bh30_80_160 <= heap_bh30_w72_13 & heap_bh30_w72_12;
      Compressor_bh30_80: Compressor_23_3
      port map ( R => CompressorOut_bh30_80_80,
                 X0 => CompressorIn_bh30_80_159,
                 X1 => CompressorIn_bh30_80_160);
   heap_bh30_w71_13 <= CompressorOut_bh30_80_80(0); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w72_14 <= CompressorOut_bh30_80_80(1); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w73_14 <= CompressorOut_bh30_80_80(2); -- cycle= 0 cp= 1.6532e-09

   CompressorIn_bh30_81_161 <= heap_bh30_w74_0 & heap_bh30_w74_12 & heap_bh30_w74_11;
   CompressorIn_bh30_81_162 <= heap_bh30_w75_13 & heap_bh30_w75_12;
      Compressor_bh30_81: Compressor_23_3
      port map ( R => CompressorOut_bh30_81_81,
                 X0 => CompressorIn_bh30_81_161,
                 X1 => CompressorIn_bh30_81_162);
   heap_bh30_w74_13 <= CompressorOut_bh30_81_81(0); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w75_14 <= CompressorOut_bh30_81_81(1); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w76_14 <= CompressorOut_bh30_81_81(2); -- cycle= 0 cp= 1.6532e-09

   CompressorIn_bh30_82_163 <= heap_bh30_w77_0 & heap_bh30_w77_12 & heap_bh30_w77_11;
   CompressorIn_bh30_82_164 <= heap_bh30_w78_13 & heap_bh30_w78_12;
      Compressor_bh30_82: Compressor_23_3
      port map ( R => CompressorOut_bh30_82_82,
                 X0 => CompressorIn_bh30_82_163,
                 X1 => CompressorIn_bh30_82_164);
   heap_bh30_w77_13 <= CompressorOut_bh30_82_82(0); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w78_14 <= CompressorOut_bh30_82_82(1); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w79_14 <= CompressorOut_bh30_82_82(2); -- cycle= 0 cp= 1.6532e-09

   CompressorIn_bh30_83_165 <= heap_bh30_w80_0 & heap_bh30_w80_12 & heap_bh30_w80_11;
   CompressorIn_bh30_83_166 <= heap_bh30_w81_13 & heap_bh30_w81_12;
      Compressor_bh30_83: Compressor_23_3
      port map ( R => CompressorOut_bh30_83_83,
                 X0 => CompressorIn_bh30_83_165,
                 X1 => CompressorIn_bh30_83_166);
   heap_bh30_w80_13 <= CompressorOut_bh30_83_83(0); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w81_14 <= CompressorOut_bh30_83_83(1); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w82_14 <= CompressorOut_bh30_83_83(2); -- cycle= 0 cp= 1.6532e-09

   CompressorIn_bh30_84_167 <= heap_bh30_w83_0 & heap_bh30_w83_12 & heap_bh30_w83_11;
   CompressorIn_bh30_84_168 <= heap_bh30_w84_13 & heap_bh30_w84_12;
      Compressor_bh30_84: Compressor_23_3
      port map ( R => CompressorOut_bh30_84_84,
                 X0 => CompressorIn_bh30_84_167,
                 X1 => CompressorIn_bh30_84_168);
   heap_bh30_w83_13 <= CompressorOut_bh30_84_84(0); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w84_14 <= CompressorOut_bh30_84_84(1); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w85_14 <= CompressorOut_bh30_84_84(2); -- cycle= 0 cp= 1.6532e-09

   CompressorIn_bh30_85_169 <= heap_bh30_w86_0 & heap_bh30_w86_12 & heap_bh30_w86_11;
   CompressorIn_bh30_85_170 <= heap_bh30_w87_13 & heap_bh30_w87_12;
      Compressor_bh30_85: Compressor_23_3
      port map ( R => CompressorOut_bh30_85_85,
                 X0 => CompressorIn_bh30_85_169,
                 X1 => CompressorIn_bh30_85_170);
   heap_bh30_w86_13 <= CompressorOut_bh30_85_85(0); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w87_14 <= CompressorOut_bh30_85_85(1); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w88_14 <= CompressorOut_bh30_85_85(2); -- cycle= 0 cp= 1.6532e-09

   CompressorIn_bh30_86_171 <= heap_bh30_w89_0 & heap_bh30_w89_12 & heap_bh30_w89_11;
   CompressorIn_bh30_86_172 <= heap_bh30_w90_12 & heap_bh30_w90_11;
      Compressor_bh30_86: Compressor_23_3
      port map ( R => CompressorOut_bh30_86_86,
                 X0 => CompressorIn_bh30_86_171,
                 X1 => CompressorIn_bh30_86_172);
   heap_bh30_w89_13 <= CompressorOut_bh30_86_86(0); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w90_13 <= CompressorOut_bh30_86_86(1); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w91_12 <= CompressorOut_bh30_86_86(2); -- cycle= 0 cp= 1.6532e-09

   CompressorIn_bh30_87_173 <= heap_bh30_w91_0 & heap_bh30_w91_11 & heap_bh30_w91_12;
   CompressorIn_bh30_87_174 <= heap_bh30_w92_0 & heap_bh30_w92_9;
      Compressor_bh30_87: Compressor_23_3
      port map ( R => CompressorOut_bh30_87_87,
                 X0 => CompressorIn_bh30_87_173,
                 X1 => CompressorIn_bh30_87_174);
   heap_bh30_w91_13 <= CompressorOut_bh30_87_87(0); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w92_10 <= CompressorOut_bh30_87_87(1); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w93_9 <= CompressorOut_bh30_87_87(2); -- cycle= 0 cp= 2.18392e-09

   CompressorIn_bh30_88_175 <= heap_bh30_w10_6 & heap_bh30_w10_5 & heap_bh30_w10_7;
   CompressorIn_bh30_88_176(0) <= heap_bh30_w11_6;
      Compressor_bh30_88: Compressor_13_3
      port map ( R => CompressorOut_bh30_88_88,
                 X0 => CompressorIn_bh30_88_175,
                 X1 => CompressorIn_bh30_88_176);
   heap_bh30_w10_8 <= CompressorOut_bh30_88_88(0); -- cycle= 0 cp= 2.16648e-09
   heap_bh30_w11_7 <= CompressorOut_bh30_88_88(1); -- cycle= 0 cp= 2.16648e-09
   heap_bh30_w12_8 <= CompressorOut_bh30_88_88(2); -- cycle= 0 cp= 2.16648e-09

   CompressorIn_bh30_89_177 <= heap_bh30_w13_6 & heap_bh30_w13_5 & heap_bh30_w13_7;
   CompressorIn_bh30_89_178(0) <= heap_bh30_w14_6;
      Compressor_bh30_89: Compressor_13_3
      port map ( R => CompressorOut_bh30_89_89,
                 X0 => CompressorIn_bh30_89_177,
                 X1 => CompressorIn_bh30_89_178);
   heap_bh30_w13_8 <= CompressorOut_bh30_89_89(0); -- cycle= 0 cp= 2.16648e-09
   heap_bh30_w14_7 <= CompressorOut_bh30_89_89(1); -- cycle= 0 cp= 2.16648e-09
   heap_bh30_w15_8 <= CompressorOut_bh30_89_89(2); -- cycle= 0 cp= 2.16648e-09

   CompressorIn_bh30_90_179 <= heap_bh30_w16_7 & heap_bh30_w16_6 & heap_bh30_w16_8;
   CompressorIn_bh30_90_180(0) <= heap_bh30_w17_7;
      Compressor_bh30_90: Compressor_13_3
      port map ( R => CompressorOut_bh30_90_90,
                 X0 => CompressorIn_bh30_90_179,
                 X1 => CompressorIn_bh30_90_180);
   heap_bh30_w16_9 <= CompressorOut_bh30_90_90(0); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w17_8 <= CompressorOut_bh30_90_90(1); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w18_9 <= CompressorOut_bh30_90_90(2); -- cycle= 0 cp= 2.18392e-09

   CompressorIn_bh30_91_181 <= heap_bh30_w19_7 & heap_bh30_w19_6 & heap_bh30_w19_8;
   CompressorIn_bh30_91_182(0) <= heap_bh30_w20_7;
      Compressor_bh30_91: Compressor_13_3
      port map ( R => CompressorOut_bh30_91_91,
                 X0 => CompressorIn_bh30_91_181,
                 X1 => CompressorIn_bh30_91_182);
   heap_bh30_w19_9 <= CompressorOut_bh30_91_91(0); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w20_8 <= CompressorOut_bh30_91_91(1); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w21_9 <= CompressorOut_bh30_91_91(2); -- cycle= 0 cp= 2.18392e-09

   CompressorIn_bh30_92_183 <= heap_bh30_w22_7 & heap_bh30_w22_6 & heap_bh30_w22_8;
   CompressorIn_bh30_92_184(0) <= heap_bh30_w23_8;
      Compressor_bh30_92: Compressor_13_3
      port map ( R => CompressorOut_bh30_92_92,
                 X0 => CompressorIn_bh30_92_183,
                 X1 => CompressorIn_bh30_92_184);
   heap_bh30_w22_9 <= CompressorOut_bh30_92_92(0); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w23_9 <= CompressorOut_bh30_92_92(1); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w24_10 <= CompressorOut_bh30_92_92(2); -- cycle= 0 cp= 2.18392e-09

   CompressorIn_bh30_93_185 <= heap_bh30_w25_8 & heap_bh30_w25_7 & heap_bh30_w25_9;
   CompressorIn_bh30_93_186(0) <= heap_bh30_w26_8;
      Compressor_bh30_93: Compressor_13_3
      port map ( R => CompressorOut_bh30_93_93,
                 X0 => CompressorIn_bh30_93_185,
                 X1 => CompressorIn_bh30_93_186);
   heap_bh30_w25_10 <= CompressorOut_bh30_93_93(0); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w26_9 <= CompressorOut_bh30_93_93(1); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w27_10 <= CompressorOut_bh30_93_93(2); -- cycle= 0 cp= 2.18392e-09

   CompressorIn_bh30_94_187 <= heap_bh30_w28_8 & heap_bh30_w28_7 & heap_bh30_w28_9;
   CompressorIn_bh30_94_188(0) <= heap_bh30_w29_8;
      Compressor_bh30_94: Compressor_13_3
      port map ( R => CompressorOut_bh30_94_94,
                 X0 => CompressorIn_bh30_94_187,
                 X1 => CompressorIn_bh30_94_188);
   heap_bh30_w28_10 <= CompressorOut_bh30_94_94(0); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w29_9 <= CompressorOut_bh30_94_94(1); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w30_10 <= CompressorOut_bh30_94_94(2); -- cycle= 0 cp= 2.18392e-09

   CompressorIn_bh30_95_189 <= heap_bh30_w31_8 & heap_bh30_w31_7 & heap_bh30_w31_9;
   CompressorIn_bh30_95_190(0) <= heap_bh30_w32_8;
      Compressor_bh30_95: Compressor_13_3
      port map ( R => CompressorOut_bh30_95_95,
                 X0 => CompressorIn_bh30_95_189,
                 X1 => CompressorIn_bh30_95_190);
   heap_bh30_w31_10 <= CompressorOut_bh30_95_95(0); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w32_9 <= CompressorOut_bh30_95_95(1); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w33_11 <= CompressorOut_bh30_95_95(2); -- cycle= 0 cp= 2.18392e-09

   CompressorIn_bh30_96_191 <= heap_bh30_w34_9 & heap_bh30_w34_8 & heap_bh30_w34_10;
   CompressorIn_bh30_96_192(0) <= heap_bh30_w35_9;
      Compressor_bh30_96: Compressor_13_3
      port map ( R => CompressorOut_bh30_96_96,
                 X0 => CompressorIn_bh30_96_191,
                 X1 => CompressorIn_bh30_96_192);
   heap_bh30_w34_11 <= CompressorOut_bh30_96_96(0); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w35_10 <= CompressorOut_bh30_96_96(1); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w36_11 <= CompressorOut_bh30_96_96(2); -- cycle= 0 cp= 2.18392e-09

   CompressorIn_bh30_97_193 <= heap_bh30_w37_9 & heap_bh30_w37_8 & heap_bh30_w37_10;
   CompressorIn_bh30_97_194(0) <= heap_bh30_w38_9;
      Compressor_bh30_97: Compressor_13_3
      port map ( R => CompressorOut_bh30_97_97,
                 X0 => CompressorIn_bh30_97_193,
                 X1 => CompressorIn_bh30_97_194);
   heap_bh30_w37_11 <= CompressorOut_bh30_97_97(0); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w38_10 <= CompressorOut_bh30_97_97(1); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w39_11 <= CompressorOut_bh30_97_97(2); -- cycle= 0 cp= 2.18392e-09

   CompressorIn_bh30_98_195 <= heap_bh30_w40_9 & heap_bh30_w40_8 & heap_bh30_w40_10;
   CompressorIn_bh30_98_196(0) <= heap_bh30_w41_9;
      Compressor_bh30_98: Compressor_13_3
      port map ( R => CompressorOut_bh30_98_98,
                 X0 => CompressorIn_bh30_98_195,
                 X1 => CompressorIn_bh30_98_196);
   heap_bh30_w40_11 <= CompressorOut_bh30_98_98(0); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w41_10 <= CompressorOut_bh30_98_98(1); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w42_11 <= CompressorOut_bh30_98_98(2); -- cycle= 0 cp= 2.18392e-09

   CompressorIn_bh30_99_197 <= heap_bh30_w43_9 & heap_bh30_w43_8 & heap_bh30_w43_10;
   CompressorIn_bh30_99_198(0) <= heap_bh30_w44_9;
      Compressor_bh30_99: Compressor_13_3
      port map ( R => CompressorOut_bh30_99_99,
                 X0 => CompressorIn_bh30_99_197,
                 X1 => CompressorIn_bh30_99_198);
   heap_bh30_w43_11 <= CompressorOut_bh30_99_99(0); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w44_10 <= CompressorOut_bh30_99_99(1); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w45_11 <= CompressorOut_bh30_99_99(2); -- cycle= 0 cp= 2.18392e-09

   CompressorIn_bh30_100_199 <= heap_bh30_w46_9 & heap_bh30_w46_8 & heap_bh30_w46_10;
   CompressorIn_bh30_100_200(0) <= heap_bh30_w47_10;
      Compressor_bh30_100: Compressor_13_3
      port map ( R => CompressorOut_bh30_100_100,
                 X0 => CompressorIn_bh30_100_199,
                 X1 => CompressorIn_bh30_100_200);
   heap_bh30_w46_11 <= CompressorOut_bh30_100_100(0); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w47_11 <= CompressorOut_bh30_100_100(1); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w48_12 <= CompressorOut_bh30_100_100(2); -- cycle= 0 cp= 2.18392e-09

   CompressorIn_bh30_101_201 <= heap_bh30_w49_10 & heap_bh30_w49_9 & heap_bh30_w49_11;
   CompressorIn_bh30_101_202(0) <= heap_bh30_w50_11;
      Compressor_bh30_101: Compressor_13_3
      port map ( R => CompressorOut_bh30_101_101,
                 X0 => CompressorIn_bh30_101_201,
                 X1 => CompressorIn_bh30_101_202);
   heap_bh30_w49_12 <= CompressorOut_bh30_101_101(0); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w50_12 <= CompressorOut_bh30_101_101(1); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w51_13 <= CompressorOut_bh30_101_101(2); -- cycle= 0 cp= 2.18392e-09

   CompressorIn_bh30_102_203 <= heap_bh30_w52_11 & heap_bh30_w52_10 & heap_bh30_w52_12;
   CompressorIn_bh30_102_204(0) <= heap_bh30_w53_11;
      Compressor_bh30_102: Compressor_13_3
      port map ( R => CompressorOut_bh30_102_102,
                 X0 => CompressorIn_bh30_102_203,
                 X1 => CompressorIn_bh30_102_204);
   heap_bh30_w52_13 <= CompressorOut_bh30_102_102(0); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w53_12 <= CompressorOut_bh30_102_102(1); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w54_13 <= CompressorOut_bh30_102_102(2); -- cycle= 0 cp= 2.18392e-09

   CompressorIn_bh30_103_205 <= heap_bh30_w55_11 & heap_bh30_w55_10 & heap_bh30_w55_12;
   CompressorIn_bh30_103_206(0) <= heap_bh30_w56_11;
      Compressor_bh30_103: Compressor_13_3
      port map ( R => CompressorOut_bh30_103_103,
                 X0 => CompressorIn_bh30_103_205,
                 X1 => CompressorIn_bh30_103_206);
   heap_bh30_w55_13 <= CompressorOut_bh30_103_103(0); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w56_12 <= CompressorOut_bh30_103_103(1); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w57_13 <= CompressorOut_bh30_103_103(2); -- cycle= 0 cp= 2.18392e-09

   CompressorIn_bh30_104_207 <= heap_bh30_w58_11 & heap_bh30_w58_10 & heap_bh30_w58_12;
   CompressorIn_bh30_104_208(0) <= heap_bh30_w59_11;
      Compressor_bh30_104: Compressor_13_3
      port map ( R => CompressorOut_bh30_104_104,
                 X0 => CompressorIn_bh30_104_207,
                 X1 => CompressorIn_bh30_104_208);
   heap_bh30_w58_13 <= CompressorOut_bh30_104_104(0); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w59_12 <= CompressorOut_bh30_104_104(1); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w60_13 <= CompressorOut_bh30_104_104(2); -- cycle= 0 cp= 2.18392e-09

   CompressorIn_bh30_105_209 <= heap_bh30_w61_11 & heap_bh30_w61_10 & heap_bh30_w61_12;
   CompressorIn_bh30_105_210(0) <= heap_bh30_w62_11;
      Compressor_bh30_105: Compressor_13_3
      port map ( R => CompressorOut_bh30_105_105,
                 X0 => CompressorIn_bh30_105_209,
                 X1 => CompressorIn_bh30_105_210);
   heap_bh30_w61_13 <= CompressorOut_bh30_105_105(0); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w62_12 <= CompressorOut_bh30_105_105(1); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w63_13 <= CompressorOut_bh30_105_105(2); -- cycle= 0 cp= 2.18392e-09

   CompressorIn_bh30_106_211 <= heap_bh30_w64_11 & heap_bh30_w64_10 & heap_bh30_w64_12;
   CompressorIn_bh30_106_212(0) <= heap_bh30_w65_11;
      Compressor_bh30_106: Compressor_13_3
      port map ( R => CompressorOut_bh30_106_106,
                 X0 => CompressorIn_bh30_106_211,
                 X1 => CompressorIn_bh30_106_212);
   heap_bh30_w64_13 <= CompressorOut_bh30_106_106(0); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w65_12 <= CompressorOut_bh30_106_106(1); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w66_13 <= CompressorOut_bh30_106_106(2); -- cycle= 0 cp= 2.18392e-09

   CompressorIn_bh30_107_213 <= heap_bh30_w67_12 & heap_bh30_w67_11 & heap_bh30_w67_13;
   CompressorIn_bh30_107_214(0) <= heap_bh30_w68_12;
      Compressor_bh30_107: Compressor_13_3
      port map ( R => CompressorOut_bh30_107_107,
                 X0 => CompressorIn_bh30_107_213,
                 X1 => CompressorIn_bh30_107_214);
   heap_bh30_w67_14 <= CompressorOut_bh30_107_107(0); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w68_13 <= CompressorOut_bh30_107_107(1); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w69_14 <= CompressorOut_bh30_107_107(2); -- cycle= 0 cp= 2.18392e-09

   CompressorIn_bh30_108_215 <= heap_bh30_w70_12 & heap_bh30_w70_11 & heap_bh30_w70_13;
   CompressorIn_bh30_108_216(0) <= heap_bh30_w71_13;
      Compressor_bh30_108: Compressor_13_3
      port map ( R => CompressorOut_bh30_108_108,
                 X0 => CompressorIn_bh30_108_215,
                 X1 => CompressorIn_bh30_108_216);
   heap_bh30_w70_14 <= CompressorOut_bh30_108_108(0); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w71_14 <= CompressorOut_bh30_108_108(1); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w72_15 <= CompressorOut_bh30_108_108(2); -- cycle= 0 cp= 2.18392e-09

   CompressorIn_bh30_109_217 <= heap_bh30_w73_13 & heap_bh30_w73_12 & heap_bh30_w73_14;
   CompressorIn_bh30_109_218(0) <= heap_bh30_w74_13;
      Compressor_bh30_109: Compressor_13_3
      port map ( R => CompressorOut_bh30_109_109,
                 X0 => CompressorIn_bh30_109_217,
                 X1 => CompressorIn_bh30_109_218);
   heap_bh30_w73_15 <= CompressorOut_bh30_109_109(0); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w74_14 <= CompressorOut_bh30_109_109(1); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w75_15 <= CompressorOut_bh30_109_109(2); -- cycle= 0 cp= 2.18392e-09

   CompressorIn_bh30_110_219 <= heap_bh30_w76_13 & heap_bh30_w76_12 & heap_bh30_w76_14;
   CompressorIn_bh30_110_220(0) <= heap_bh30_w77_13;
      Compressor_bh30_110: Compressor_13_3
      port map ( R => CompressorOut_bh30_110_110,
                 X0 => CompressorIn_bh30_110_219,
                 X1 => CompressorIn_bh30_110_220);
   heap_bh30_w76_15 <= CompressorOut_bh30_110_110(0); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w77_14 <= CompressorOut_bh30_110_110(1); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w78_15 <= CompressorOut_bh30_110_110(2); -- cycle= 0 cp= 2.18392e-09

   CompressorIn_bh30_111_221 <= heap_bh30_w79_13 & heap_bh30_w79_12 & heap_bh30_w79_14;
   CompressorIn_bh30_111_222(0) <= heap_bh30_w80_13;
      Compressor_bh30_111: Compressor_13_3
      port map ( R => CompressorOut_bh30_111_111,
                 X0 => CompressorIn_bh30_111_221,
                 X1 => CompressorIn_bh30_111_222);
   heap_bh30_w79_15 <= CompressorOut_bh30_111_111(0); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w80_14 <= CompressorOut_bh30_111_111(1); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w81_15 <= CompressorOut_bh30_111_111(2); -- cycle= 0 cp= 2.18392e-09

   CompressorIn_bh30_112_223 <= heap_bh30_w82_13 & heap_bh30_w82_12 & heap_bh30_w82_14;
   CompressorIn_bh30_112_224(0) <= heap_bh30_w83_13;
      Compressor_bh30_112: Compressor_13_3
      port map ( R => CompressorOut_bh30_112_112,
                 X0 => CompressorIn_bh30_112_223,
                 X1 => CompressorIn_bh30_112_224);
   heap_bh30_w82_15 <= CompressorOut_bh30_112_112(0); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w83_14 <= CompressorOut_bh30_112_112(1); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w84_15 <= CompressorOut_bh30_112_112(2); -- cycle= 0 cp= 2.18392e-09

   CompressorIn_bh30_113_225 <= heap_bh30_w85_13 & heap_bh30_w85_12 & heap_bh30_w85_14;
   CompressorIn_bh30_113_226(0) <= heap_bh30_w86_13;
      Compressor_bh30_113: Compressor_13_3
      port map ( R => CompressorOut_bh30_113_113,
                 X0 => CompressorIn_bh30_113_225,
                 X1 => CompressorIn_bh30_113_226);
   heap_bh30_w85_15 <= CompressorOut_bh30_113_113(0); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w86_14 <= CompressorOut_bh30_113_113(1); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w87_15 <= CompressorOut_bh30_113_113(2); -- cycle= 0 cp= 2.18392e-09

   CompressorIn_bh30_114_227 <= heap_bh30_w88_13 & heap_bh30_w88_12 & heap_bh30_w88_14;
   CompressorIn_bh30_114_228(0) <= heap_bh30_w89_13;
      Compressor_bh30_114: Compressor_13_3
      port map ( R => CompressorOut_bh30_114_114,
                 X0 => CompressorIn_bh30_114_227,
                 X1 => CompressorIn_bh30_114_228);
   heap_bh30_w88_15 <= CompressorOut_bh30_114_114(0); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w89_14 <= CompressorOut_bh30_114_114(1); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w90_14 <= CompressorOut_bh30_114_114(2); -- cycle= 0 cp= 2.18392e-09

   CompressorIn_bh30_115_229 <= heap_bh30_w33_10 & heap_bh30_w33_11 & heap_bh30_w33_7 & heap_bh30_w33_6 & heap_bh30_w33_5 & heap_bh30_w33_4;
      Compressor_bh30_115: Compressor_6_3
      port map ( R => CompressorOut_bh30_115_115,
                 X0 => CompressorIn_bh30_115_229);
   heap_bh30_w33_12 <= CompressorOut_bh30_115_115(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w34_12 <= CompressorOut_bh30_115_115(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w35_11 <= CompressorOut_bh30_115_115(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_116_230 <= heap_bh30_w36_10 & heap_bh30_w36_11 & heap_bh30_w36_7 & heap_bh30_w36_6 & heap_bh30_w36_5 & heap_bh30_w36_4;
      Compressor_bh30_116: Compressor_6_3
      port map ( R => CompressorOut_bh30_116_116,
                 X0 => CompressorIn_bh30_116_230);
   heap_bh30_w36_12 <= CompressorOut_bh30_116_116(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w37_12 <= CompressorOut_bh30_116_116(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w38_11 <= CompressorOut_bh30_116_116(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_117_231 <= heap_bh30_w39_10 & heap_bh30_w39_11 & heap_bh30_w39_7 & heap_bh30_w39_6 & heap_bh30_w39_5 & heap_bh30_w39_4;
      Compressor_bh30_117: Compressor_6_3
      port map ( R => CompressorOut_bh30_117_117,
                 X0 => CompressorIn_bh30_117_231);
   heap_bh30_w39_12 <= CompressorOut_bh30_117_117(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w40_12 <= CompressorOut_bh30_117_117(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w41_11 <= CompressorOut_bh30_117_117(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_118_232 <= heap_bh30_w42_10 & heap_bh30_w42_11 & heap_bh30_w42_7 & heap_bh30_w42_6 & heap_bh30_w42_5 & heap_bh30_w42_4;
      Compressor_bh30_118: Compressor_6_3
      port map ( R => CompressorOut_bh30_118_118,
                 X0 => CompressorIn_bh30_118_232);
   heap_bh30_w42_12 <= CompressorOut_bh30_118_118(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w43_12 <= CompressorOut_bh30_118_118(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w44_11 <= CompressorOut_bh30_118_118(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_119_233 <= heap_bh30_w45_10 & heap_bh30_w45_11 & heap_bh30_w45_7 & heap_bh30_w45_6 & heap_bh30_w45_5 & heap_bh30_w45_4;
      Compressor_bh30_119: Compressor_6_3
      port map ( R => CompressorOut_bh30_119_119,
                 X0 => CompressorIn_bh30_119_233);
   heap_bh30_w45_12 <= CompressorOut_bh30_119_119(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w46_12 <= CompressorOut_bh30_119_119(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w47_12 <= CompressorOut_bh30_119_119(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_120_234 <= heap_bh30_w47_11 & heap_bh30_w47_7 & heap_bh30_w47_6 & heap_bh30_w47_5 & heap_bh30_w47_4 & heap_bh30_w47_3;
      Compressor_bh30_120: Compressor_6_3
      port map ( R => CompressorOut_bh30_120_120,
                 X0 => CompressorIn_bh30_120_234);
   heap_bh30_w47_13 <= CompressorOut_bh30_120_120(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w48_13 <= CompressorOut_bh30_120_120(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w49_13 <= CompressorOut_bh30_120_120(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_121_235 <= heap_bh30_w48_11 & heap_bh30_w48_12 & heap_bh30_w48_8 & heap_bh30_w48_7 & heap_bh30_w48_6 & heap_bh30_w48_5;
      Compressor_bh30_121: Compressor_6_3
      port map ( R => CompressorOut_bh30_121_121,
                 X0 => CompressorIn_bh30_121_235);
   heap_bh30_w48_14 <= CompressorOut_bh30_121_121(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w49_14 <= CompressorOut_bh30_121_121(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w50_13 <= CompressorOut_bh30_121_121(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_122_236 <= heap_bh30_w49_12 & heap_bh30_w49_8 & heap_bh30_w49_7 & heap_bh30_w49_6 & heap_bh30_w49_5 & heap_bh30_w49_4;
      Compressor_bh30_122: Compressor_6_3
      port map ( R => CompressorOut_bh30_122_122,
                 X0 => CompressorIn_bh30_122_236);
   heap_bh30_w49_15 <= CompressorOut_bh30_122_122(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w50_14 <= CompressorOut_bh30_122_122(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w51_14 <= CompressorOut_bh30_122_122(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_123_237 <= heap_bh30_w50_12 & heap_bh30_w50_8 & heap_bh30_w50_7 & heap_bh30_w50_6 & heap_bh30_w50_5 & heap_bh30_w50_4;
      Compressor_bh30_123: Compressor_6_3
      port map ( R => CompressorOut_bh30_123_123,
                 X0 => CompressorIn_bh30_123_237);
   heap_bh30_w50_15 <= CompressorOut_bh30_123_123(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w51_15 <= CompressorOut_bh30_123_123(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w52_14 <= CompressorOut_bh30_123_123(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_124_238 <= heap_bh30_w51_12 & heap_bh30_w51_13 & heap_bh30_w51_9 & heap_bh30_w51_8 & heap_bh30_w51_7 & heap_bh30_w51_6;
      Compressor_bh30_124: Compressor_6_3
      port map ( R => CompressorOut_bh30_124_124,
                 X0 => CompressorIn_bh30_124_238);
   heap_bh30_w51_16 <= CompressorOut_bh30_124_124(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w52_15 <= CompressorOut_bh30_124_124(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w53_13 <= CompressorOut_bh30_124_124(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_125_239 <= heap_bh30_w52_13 & heap_bh30_w52_9 & heap_bh30_w52_8 & heap_bh30_w52_7 & heap_bh30_w52_6 & heap_bh30_w52_5;
      Compressor_bh30_125: Compressor_6_3
      port map ( R => CompressorOut_bh30_125_125,
                 X0 => CompressorIn_bh30_125_239);
   heap_bh30_w52_16 <= CompressorOut_bh30_125_125(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w53_14 <= CompressorOut_bh30_125_125(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w54_14 <= CompressorOut_bh30_125_125(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_126_240 <= heap_bh30_w53_12 & heap_bh30_w53_8 & heap_bh30_w53_7 & heap_bh30_w53_6 & heap_bh30_w53_5 & heap_bh30_w53_4;
      Compressor_bh30_126: Compressor_6_3
      port map ( R => CompressorOut_bh30_126_126,
                 X0 => CompressorIn_bh30_126_240);
   heap_bh30_w53_15 <= CompressorOut_bh30_126_126(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w54_15 <= CompressorOut_bh30_126_126(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w55_14 <= CompressorOut_bh30_126_126(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_127_241 <= heap_bh30_w54_12 & heap_bh30_w54_13 & heap_bh30_w54_9 & heap_bh30_w54_8 & heap_bh30_w54_7 & heap_bh30_w54_6;
      Compressor_bh30_127: Compressor_6_3
      port map ( R => CompressorOut_bh30_127_127,
                 X0 => CompressorIn_bh30_127_241);
   heap_bh30_w54_16 <= CompressorOut_bh30_127_127(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w55_15 <= CompressorOut_bh30_127_127(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w56_13 <= CompressorOut_bh30_127_127(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_128_242 <= heap_bh30_w55_13 & heap_bh30_w55_9 & heap_bh30_w55_8 & heap_bh30_w55_7 & heap_bh30_w55_6 & heap_bh30_w55_5;
      Compressor_bh30_128: Compressor_6_3
      port map ( R => CompressorOut_bh30_128_128,
                 X0 => CompressorIn_bh30_128_242);
   heap_bh30_w55_16 <= CompressorOut_bh30_128_128(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w56_14 <= CompressorOut_bh30_128_128(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w57_14 <= CompressorOut_bh30_128_128(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_129_243 <= heap_bh30_w56_12 & heap_bh30_w56_8 & heap_bh30_w56_7 & heap_bh30_w56_6 & heap_bh30_w56_5 & heap_bh30_w56_4;
      Compressor_bh30_129: Compressor_6_3
      port map ( R => CompressorOut_bh30_129_129,
                 X0 => CompressorIn_bh30_129_243);
   heap_bh30_w56_15 <= CompressorOut_bh30_129_129(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w57_15 <= CompressorOut_bh30_129_129(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w58_14 <= CompressorOut_bh30_129_129(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_130_244 <= heap_bh30_w57_12 & heap_bh30_w57_13 & heap_bh30_w57_9 & heap_bh30_w57_8 & heap_bh30_w57_7 & heap_bh30_w57_6;
      Compressor_bh30_130: Compressor_6_3
      port map ( R => CompressorOut_bh30_130_130,
                 X0 => CompressorIn_bh30_130_244);
   heap_bh30_w57_16 <= CompressorOut_bh30_130_130(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w58_15 <= CompressorOut_bh30_130_130(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w59_13 <= CompressorOut_bh30_130_130(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_131_245 <= heap_bh30_w58_13 & heap_bh30_w58_9 & heap_bh30_w58_8 & heap_bh30_w58_7 & heap_bh30_w58_6 & heap_bh30_w58_5;
      Compressor_bh30_131: Compressor_6_3
      port map ( R => CompressorOut_bh30_131_131,
                 X0 => CompressorIn_bh30_131_245);
   heap_bh30_w58_16 <= CompressorOut_bh30_131_131(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w59_14 <= CompressorOut_bh30_131_131(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w60_14 <= CompressorOut_bh30_131_131(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_132_246 <= heap_bh30_w59_12 & heap_bh30_w59_8 & heap_bh30_w59_7 & heap_bh30_w59_6 & heap_bh30_w59_5 & heap_bh30_w59_4;
      Compressor_bh30_132: Compressor_6_3
      port map ( R => CompressorOut_bh30_132_132,
                 X0 => CompressorIn_bh30_132_246);
   heap_bh30_w59_15 <= CompressorOut_bh30_132_132(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w60_15 <= CompressorOut_bh30_132_132(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w61_14 <= CompressorOut_bh30_132_132(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_133_247 <= heap_bh30_w60_12 & heap_bh30_w60_13 & heap_bh30_w60_9 & heap_bh30_w60_8 & heap_bh30_w60_7 & heap_bh30_w60_6;
      Compressor_bh30_133: Compressor_6_3
      port map ( R => CompressorOut_bh30_133_133,
                 X0 => CompressorIn_bh30_133_247);
   heap_bh30_w60_16 <= CompressorOut_bh30_133_133(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w61_15 <= CompressorOut_bh30_133_133(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w62_13 <= CompressorOut_bh30_133_133(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_134_248 <= heap_bh30_w61_13 & heap_bh30_w61_9 & heap_bh30_w61_8 & heap_bh30_w61_7 & heap_bh30_w61_6 & heap_bh30_w61_5;
      Compressor_bh30_134: Compressor_6_3
      port map ( R => CompressorOut_bh30_134_134,
                 X0 => CompressorIn_bh30_134_248);
   heap_bh30_w61_16 <= CompressorOut_bh30_134_134(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w62_14 <= CompressorOut_bh30_134_134(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w63_14 <= CompressorOut_bh30_134_134(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_135_249 <= heap_bh30_w62_12 & heap_bh30_w62_8 & heap_bh30_w62_7 & heap_bh30_w62_6 & heap_bh30_w62_5 & heap_bh30_w62_4;
      Compressor_bh30_135: Compressor_6_3
      port map ( R => CompressorOut_bh30_135_135,
                 X0 => CompressorIn_bh30_135_249);
   heap_bh30_w62_15 <= CompressorOut_bh30_135_135(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w63_15 <= CompressorOut_bh30_135_135(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w64_14 <= CompressorOut_bh30_135_135(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_136_250 <= heap_bh30_w63_12 & heap_bh30_w63_13 & heap_bh30_w63_9 & heap_bh30_w63_8 & heap_bh30_w63_7 & heap_bh30_w63_6;
      Compressor_bh30_136: Compressor_6_3
      port map ( R => CompressorOut_bh30_136_136,
                 X0 => CompressorIn_bh30_136_250);
   heap_bh30_w63_16 <= CompressorOut_bh30_136_136(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w64_15 <= CompressorOut_bh30_136_136(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w65_13 <= CompressorOut_bh30_136_136(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_137_251 <= heap_bh30_w64_13 & heap_bh30_w64_9 & heap_bh30_w64_8 & heap_bh30_w64_7 & heap_bh30_w64_6 & heap_bh30_w64_5;
      Compressor_bh30_137: Compressor_6_3
      port map ( R => CompressorOut_bh30_137_137,
                 X0 => CompressorIn_bh30_137_251);
   heap_bh30_w64_16 <= CompressorOut_bh30_137_137(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w65_14 <= CompressorOut_bh30_137_137(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w66_14 <= CompressorOut_bh30_137_137(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_138_252 <= heap_bh30_w65_12 & heap_bh30_w65_8 & heap_bh30_w65_7 & heap_bh30_w65_6 & heap_bh30_w65_5 & heap_bh30_w65_4;
      Compressor_bh30_138: Compressor_6_3
      port map ( R => CompressorOut_bh30_138_138,
                 X0 => CompressorIn_bh30_138_252);
   heap_bh30_w65_15 <= CompressorOut_bh30_138_138(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w66_15 <= CompressorOut_bh30_138_138(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w67_15 <= CompressorOut_bh30_138_138(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_139_253 <= heap_bh30_w66_12 & heap_bh30_w66_13 & heap_bh30_w66_9 & heap_bh30_w66_8 & heap_bh30_w66_7 & heap_bh30_w66_6;
      Compressor_bh30_139: Compressor_6_3
      port map ( R => CompressorOut_bh30_139_139,
                 X0 => CompressorIn_bh30_139_253);
   heap_bh30_w66_16 <= CompressorOut_bh30_139_139(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w67_16 <= CompressorOut_bh30_139_139(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w68_14 <= CompressorOut_bh30_139_139(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_140_254 <= heap_bh30_w67_14 & heap_bh30_w67_10 & heap_bh30_w67_9 & heap_bh30_w67_8 & heap_bh30_w67_7 & heap_bh30_w67_6;
      Compressor_bh30_140: Compressor_6_3
      port map ( R => CompressorOut_bh30_140_140,
                 X0 => CompressorIn_bh30_140_254);
   heap_bh30_w67_17 <= CompressorOut_bh30_140_140(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w68_15 <= CompressorOut_bh30_140_140(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w69_15 <= CompressorOut_bh30_140_140(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_141_255 <= heap_bh30_w68_13 & heap_bh30_w68_9 & heap_bh30_w68_8 & heap_bh30_w68_7 & heap_bh30_w68_6 & heap_bh30_w68_5;
      Compressor_bh30_141: Compressor_6_3
      port map ( R => CompressorOut_bh30_141_141,
                 X0 => CompressorIn_bh30_141_255);
   heap_bh30_w68_16 <= CompressorOut_bh30_141_141(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w69_16 <= CompressorOut_bh30_141_141(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w70_15 <= CompressorOut_bh30_141_141(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_142_256 <= heap_bh30_w69_13 & heap_bh30_w69_14 & heap_bh30_w69_10 & heap_bh30_w69_9 & heap_bh30_w69_8 & heap_bh30_w69_7;
      Compressor_bh30_142: Compressor_6_3
      port map ( R => CompressorOut_bh30_142_142,
                 X0 => CompressorIn_bh30_142_256);
   heap_bh30_w69_17 <= CompressorOut_bh30_142_142(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w70_16 <= CompressorOut_bh30_142_142(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w71_15 <= CompressorOut_bh30_142_142(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_143_257 <= heap_bh30_w70_14 & heap_bh30_w70_10 & heap_bh30_w70_9 & heap_bh30_w70_8 & heap_bh30_w70_7 & heap_bh30_w70_6;
      Compressor_bh30_143: Compressor_6_3
      port map ( R => CompressorOut_bh30_143_143,
                 X0 => CompressorIn_bh30_143_257);
   heap_bh30_w70_17 <= CompressorOut_bh30_143_143(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w71_16 <= CompressorOut_bh30_143_143(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w72_16 <= CompressorOut_bh30_143_143(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_144_258 <= heap_bh30_w71_14 & heap_bh30_w71_10 & heap_bh30_w71_9 & heap_bh30_w71_8 & heap_bh30_w71_7 & heap_bh30_w71_6;
      Compressor_bh30_144: Compressor_6_3
      port map ( R => CompressorOut_bh30_144_144,
                 X0 => CompressorIn_bh30_144_258);
   heap_bh30_w71_17 <= CompressorOut_bh30_144_144(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w72_17 <= CompressorOut_bh30_144_144(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w73_16 <= CompressorOut_bh30_144_144(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_145_259 <= heap_bh30_w72_14 & heap_bh30_w72_15 & heap_bh30_w72_11 & heap_bh30_w72_10 & heap_bh30_w72_9 & heap_bh30_w72_8;
      Compressor_bh30_145: Compressor_6_3
      port map ( R => CompressorOut_bh30_145_145,
                 X0 => CompressorIn_bh30_145_259);
   heap_bh30_w72_18 <= CompressorOut_bh30_145_145(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w73_17 <= CompressorOut_bh30_145_145(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w74_15 <= CompressorOut_bh30_145_145(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_146_260 <= heap_bh30_w73_15 & heap_bh30_w73_11 & heap_bh30_w73_10 & heap_bh30_w73_9 & heap_bh30_w73_8 & heap_bh30_w73_7;
      Compressor_bh30_146: Compressor_6_3
      port map ( R => CompressorOut_bh30_146_146,
                 X0 => CompressorIn_bh30_146_260);
   heap_bh30_w73_18 <= CompressorOut_bh30_146_146(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w74_16 <= CompressorOut_bh30_146_146(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w75_16 <= CompressorOut_bh30_146_146(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_147_261 <= heap_bh30_w74_14 & heap_bh30_w74_10 & heap_bh30_w74_9 & heap_bh30_w74_8 & heap_bh30_w74_7 & heap_bh30_w74_6;
      Compressor_bh30_147: Compressor_6_3
      port map ( R => CompressorOut_bh30_147_147,
                 X0 => CompressorIn_bh30_147_261);
   heap_bh30_w74_17 <= CompressorOut_bh30_147_147(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w75_17 <= CompressorOut_bh30_147_147(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w76_16 <= CompressorOut_bh30_147_147(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_148_262 <= heap_bh30_w75_14 & heap_bh30_w75_15 & heap_bh30_w75_11 & heap_bh30_w75_10 & heap_bh30_w75_9 & heap_bh30_w75_8;
      Compressor_bh30_148: Compressor_6_3
      port map ( R => CompressorOut_bh30_148_148,
                 X0 => CompressorIn_bh30_148_262);
   heap_bh30_w75_18 <= CompressorOut_bh30_148_148(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w76_17 <= CompressorOut_bh30_148_148(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w77_15 <= CompressorOut_bh30_148_148(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_149_263 <= heap_bh30_w76_15 & heap_bh30_w76_11 & heap_bh30_w76_10 & heap_bh30_w76_9 & heap_bh30_w76_8 & heap_bh30_w76_7;
      Compressor_bh30_149: Compressor_6_3
      port map ( R => CompressorOut_bh30_149_149,
                 X0 => CompressorIn_bh30_149_263);
   heap_bh30_w76_18 <= CompressorOut_bh30_149_149(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w77_16 <= CompressorOut_bh30_149_149(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w78_16 <= CompressorOut_bh30_149_149(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_150_264 <= heap_bh30_w77_14 & heap_bh30_w77_10 & heap_bh30_w77_9 & heap_bh30_w77_8 & heap_bh30_w77_7 & heap_bh30_w77_6;
      Compressor_bh30_150: Compressor_6_3
      port map ( R => CompressorOut_bh30_150_150,
                 X0 => CompressorIn_bh30_150_264);
   heap_bh30_w77_17 <= CompressorOut_bh30_150_150(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w78_17 <= CompressorOut_bh30_150_150(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w79_16 <= CompressorOut_bh30_150_150(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_151_265 <= heap_bh30_w78_14 & heap_bh30_w78_15 & heap_bh30_w78_11 & heap_bh30_w78_10 & heap_bh30_w78_9 & heap_bh30_w78_8;
      Compressor_bh30_151: Compressor_6_3
      port map ( R => CompressorOut_bh30_151_151,
                 X0 => CompressorIn_bh30_151_265);
   heap_bh30_w78_18 <= CompressorOut_bh30_151_151(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w79_17 <= CompressorOut_bh30_151_151(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w80_15 <= CompressorOut_bh30_151_151(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_152_266 <= heap_bh30_w79_15 & heap_bh30_w79_11 & heap_bh30_w79_10 & heap_bh30_w79_9 & heap_bh30_w79_8 & heap_bh30_w79_7;
      Compressor_bh30_152: Compressor_6_3
      port map ( R => CompressorOut_bh30_152_152,
                 X0 => CompressorIn_bh30_152_266);
   heap_bh30_w79_18 <= CompressorOut_bh30_152_152(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w80_16 <= CompressorOut_bh30_152_152(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w81_16 <= CompressorOut_bh30_152_152(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_153_267 <= heap_bh30_w80_14 & heap_bh30_w80_10 & heap_bh30_w80_9 & heap_bh30_w80_8 & heap_bh30_w80_7 & heap_bh30_w80_6;
      Compressor_bh30_153: Compressor_6_3
      port map ( R => CompressorOut_bh30_153_153,
                 X0 => CompressorIn_bh30_153_267);
   heap_bh30_w80_17 <= CompressorOut_bh30_153_153(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w81_17 <= CompressorOut_bh30_153_153(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w82_16 <= CompressorOut_bh30_153_153(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_154_268 <= heap_bh30_w81_14 & heap_bh30_w81_15 & heap_bh30_w81_11 & heap_bh30_w81_10 & heap_bh30_w81_9 & heap_bh30_w81_8;
      Compressor_bh30_154: Compressor_6_3
      port map ( R => CompressorOut_bh30_154_154,
                 X0 => CompressorIn_bh30_154_268);
   heap_bh30_w81_18 <= CompressorOut_bh30_154_154(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w82_17 <= CompressorOut_bh30_154_154(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w83_15 <= CompressorOut_bh30_154_154(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_155_269 <= heap_bh30_w82_15 & heap_bh30_w82_11 & heap_bh30_w82_10 & heap_bh30_w82_9 & heap_bh30_w82_8 & heap_bh30_w82_7;
      Compressor_bh30_155: Compressor_6_3
      port map ( R => CompressorOut_bh30_155_155,
                 X0 => CompressorIn_bh30_155_269);
   heap_bh30_w82_18 <= CompressorOut_bh30_155_155(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w83_16 <= CompressorOut_bh30_155_155(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w84_16 <= CompressorOut_bh30_155_155(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_156_270 <= heap_bh30_w83_14 & heap_bh30_w83_10 & heap_bh30_w83_9 & heap_bh30_w83_8 & heap_bh30_w83_7 & heap_bh30_w83_6;
      Compressor_bh30_156: Compressor_6_3
      port map ( R => CompressorOut_bh30_156_156,
                 X0 => CompressorIn_bh30_156_270);
   heap_bh30_w83_17 <= CompressorOut_bh30_156_156(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w84_17 <= CompressorOut_bh30_156_156(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w85_16 <= CompressorOut_bh30_156_156(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_157_271 <= heap_bh30_w84_14 & heap_bh30_w84_15 & heap_bh30_w84_11 & heap_bh30_w84_10 & heap_bh30_w84_9 & heap_bh30_w84_8;
      Compressor_bh30_157: Compressor_6_3
      port map ( R => CompressorOut_bh30_157_157,
                 X0 => CompressorIn_bh30_157_271);
   heap_bh30_w84_18 <= CompressorOut_bh30_157_157(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w85_17 <= CompressorOut_bh30_157_157(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w86_15 <= CompressorOut_bh30_157_157(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_158_272 <= heap_bh30_w85_15 & heap_bh30_w85_11 & heap_bh30_w85_10 & heap_bh30_w85_9 & heap_bh30_w85_8 & heap_bh30_w85_7;
      Compressor_bh30_158: Compressor_6_3
      port map ( R => CompressorOut_bh30_158_158,
                 X0 => CompressorIn_bh30_158_272);
   heap_bh30_w85_18 <= CompressorOut_bh30_158_158(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w86_16 <= CompressorOut_bh30_158_158(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w87_16 <= CompressorOut_bh30_158_158(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_159_273 <= heap_bh30_w86_14 & heap_bh30_w86_10 & heap_bh30_w86_9 & heap_bh30_w86_8 & heap_bh30_w86_7 & heap_bh30_w86_6;
      Compressor_bh30_159: Compressor_6_3
      port map ( R => CompressorOut_bh30_159_159,
                 X0 => CompressorIn_bh30_159_273);
   heap_bh30_w86_17 <= CompressorOut_bh30_159_159(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w87_17 <= CompressorOut_bh30_159_159(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w88_16 <= CompressorOut_bh30_159_159(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_160_274 <= heap_bh30_w87_14 & heap_bh30_w87_15 & heap_bh30_w87_11 & heap_bh30_w87_10 & heap_bh30_w87_9 & heap_bh30_w87_8;
      Compressor_bh30_160: Compressor_6_3
      port map ( R => CompressorOut_bh30_160_160,
                 X0 => CompressorIn_bh30_160_274);
   heap_bh30_w87_18 <= CompressorOut_bh30_160_160(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w88_17 <= CompressorOut_bh30_160_160(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w89_15 <= CompressorOut_bh30_160_160(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_161_275 <= heap_bh30_w88_15 & heap_bh30_w88_11 & heap_bh30_w88_10 & heap_bh30_w88_9 & heap_bh30_w88_8 & heap_bh30_w88_7;
      Compressor_bh30_161: Compressor_6_3
      port map ( R => CompressorOut_bh30_161_161,
                 X0 => CompressorIn_bh30_161_275);
   heap_bh30_w88_18 <= CompressorOut_bh30_161_161(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w89_16 <= CompressorOut_bh30_161_161(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w90_15 <= CompressorOut_bh30_161_161(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_162_276 <= heap_bh30_w89_14 & heap_bh30_w89_10 & heap_bh30_w89_9 & heap_bh30_w89_8 & heap_bh30_w89_7 & heap_bh30_w89_6;
      Compressor_bh30_162: Compressor_6_3
      port map ( R => CompressorOut_bh30_162_162,
                 X0 => CompressorIn_bh30_162_276);
   heap_bh30_w89_17 <= CompressorOut_bh30_162_162(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w90_16 <= CompressorOut_bh30_162_162(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w91_14 <= CompressorOut_bh30_162_162(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_163_277 <= heap_bh30_w90_13 & heap_bh30_w90_14 & heap_bh30_w90_10 & heap_bh30_w90_9 & heap_bh30_w90_8 & heap_bh30_w90_7;
      Compressor_bh30_163: Compressor_6_3
      port map ( R => CompressorOut_bh30_163_163,
                 X0 => CompressorIn_bh30_163_277);
   heap_bh30_w90_17 <= CompressorOut_bh30_163_163(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w91_15 <= CompressorOut_bh30_163_163(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w92_11 <= CompressorOut_bh30_163_163(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_164_278 <= heap_bh30_w91_13 & heap_bh30_w91_10 & heap_bh30_w91_9 & heap_bh30_w91_8 & heap_bh30_w91_7 & heap_bh30_w91_6;
      Compressor_bh30_164: Compressor_6_3
      port map ( R => CompressorOut_bh30_164_164,
                 X0 => CompressorIn_bh30_164_278);
   heap_bh30_w91_16 <= CompressorOut_bh30_164_164(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w92_12 <= CompressorOut_bh30_164_164(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w93_10 <= CompressorOut_bh30_164_164(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_165_279 <= heap_bh30_w92_10 & heap_bh30_w92_8 & heap_bh30_w92_7 & heap_bh30_w92_6 & heap_bh30_w92_5 & heap_bh30_w92_4;
      Compressor_bh30_165: Compressor_6_3
      port map ( R => CompressorOut_bh30_165_165,
                 X0 => CompressorIn_bh30_165_279);
   heap_bh30_w92_13 <= CompressorOut_bh30_165_165(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w93_11 <= CompressorOut_bh30_165_165(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w94_9 <= CompressorOut_bh30_165_165(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_166_280 <= heap_bh30_w93_0 & heap_bh30_w93_9 & heap_bh30_w93_8 & heap_bh30_w93_7 & heap_bh30_w93_6 & heap_bh30_w93_5;
      Compressor_bh30_166: Compressor_6_3
      port map ( R => CompressorOut_bh30_166_166,
                 X0 => CompressorIn_bh30_166_280);
   heap_bh30_w93_12 <= CompressorOut_bh30_166_166(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w94_10 <= CompressorOut_bh30_166_166(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w95_8 <= CompressorOut_bh30_166_166(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_167_281 <= heap_bh30_w94_0 & heap_bh30_w94_8 & heap_bh30_w94_7 & heap_bh30_w94_6 & heap_bh30_w94_5 & heap_bh30_w94_4;
      Compressor_bh30_167: Compressor_6_3
      port map ( R => CompressorOut_bh30_167_167,
                 X0 => CompressorIn_bh30_167_281);
   heap_bh30_w94_11 <= CompressorOut_bh30_167_167(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w95_9 <= CompressorOut_bh30_167_167(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w96_8 <= CompressorOut_bh30_167_167(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_168_282 <= heap_bh30_w95_7 & heap_bh30_w95_6 & heap_bh30_w95_5 & heap_bh30_w95_4 & heap_bh30_w95_3 & heap_bh30_w95_2;
      Compressor_bh30_168: Compressor_6_3
      port map ( R => CompressorOut_bh30_168_168,
                 X0 => CompressorIn_bh30_168_282);
   heap_bh30_w95_10 <= CompressorOut_bh30_168_168(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w96_9 <= CompressorOut_bh30_168_168(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w97_8 <= CompressorOut_bh30_168_168(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_169_283 <= heap_bh30_w96_7 & heap_bh30_w96_6 & heap_bh30_w96_5 & heap_bh30_w96_4 & heap_bh30_w96_3 & heap_bh30_w96_2;
      Compressor_bh30_169: Compressor_6_3
      port map ( R => CompressorOut_bh30_169_169,
                 X0 => CompressorIn_bh30_169_283);
   heap_bh30_w96_10 <= CompressorOut_bh30_169_169(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w97_9 <= CompressorOut_bh30_169_169(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w98_8 <= CompressorOut_bh30_169_169(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_170_284 <= heap_bh30_w97_7 & heap_bh30_w97_6 & heap_bh30_w97_5 & heap_bh30_w97_4 & heap_bh30_w97_3 & heap_bh30_w97_2;
      Compressor_bh30_170: Compressor_6_3
      port map ( R => CompressorOut_bh30_170_170,
                 X0 => CompressorIn_bh30_170_284);
   heap_bh30_w97_10 <= CompressorOut_bh30_170_170(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w98_9 <= CompressorOut_bh30_170_170(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w99_8 <= CompressorOut_bh30_170_170(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_171_285 <= heap_bh30_w98_7 & heap_bh30_w98_6 & heap_bh30_w98_5 & heap_bh30_w98_4 & heap_bh30_w98_3 & heap_bh30_w98_2;
      Compressor_bh30_171: Compressor_6_3
      port map ( R => CompressorOut_bh30_171_171,
                 X0 => CompressorIn_bh30_171_285);
   heap_bh30_w98_10 <= CompressorOut_bh30_171_171(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w99_9 <= CompressorOut_bh30_171_171(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w100_8 <= CompressorOut_bh30_171_171(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_172_286 <= heap_bh30_w99_7 & heap_bh30_w99_6 & heap_bh30_w99_5 & heap_bh30_w99_4 & heap_bh30_w99_3 & heap_bh30_w99_2;
      Compressor_bh30_172: Compressor_6_3
      port map ( R => CompressorOut_bh30_172_172,
                 X0 => CompressorIn_bh30_172_286);
   heap_bh30_w99_10 <= CompressorOut_bh30_172_172(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w100_9 <= CompressorOut_bh30_172_172(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w101_8 <= CompressorOut_bh30_172_172(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_173_287 <= heap_bh30_w100_7 & heap_bh30_w100_6 & heap_bh30_w100_5 & heap_bh30_w100_4 & heap_bh30_w100_3 & heap_bh30_w100_2;
      Compressor_bh30_173: Compressor_6_3
      port map ( R => CompressorOut_bh30_173_173,
                 X0 => CompressorIn_bh30_173_287);
   heap_bh30_w100_10 <= CompressorOut_bh30_173_173(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w101_9 <= CompressorOut_bh30_173_173(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w102_8 <= CompressorOut_bh30_173_173(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_174_288 <= heap_bh30_w101_7 & heap_bh30_w101_6 & heap_bh30_w101_5 & heap_bh30_w101_4 & heap_bh30_w101_3 & heap_bh30_w101_2;
      Compressor_bh30_174: Compressor_6_3
      port map ( R => CompressorOut_bh30_174_174,
                 X0 => CompressorIn_bh30_174_288);
   heap_bh30_w101_10 <= CompressorOut_bh30_174_174(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w102_9 <= CompressorOut_bh30_174_174(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w103_8 <= CompressorOut_bh30_174_174(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_175_289 <= heap_bh30_w102_7 & heap_bh30_w102_6 & heap_bh30_w102_5 & heap_bh30_w102_4 & heap_bh30_w102_3 & heap_bh30_w102_2;
      Compressor_bh30_175: Compressor_6_3
      port map ( R => CompressorOut_bh30_175_175,
                 X0 => CompressorIn_bh30_175_289);
   heap_bh30_w102_10 <= CompressorOut_bh30_175_175(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w103_9 <= CompressorOut_bh30_175_175(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w104_8 <= CompressorOut_bh30_175_175(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_176_290 <= heap_bh30_w103_7 & heap_bh30_w103_6 & heap_bh30_w103_5 & heap_bh30_w103_4 & heap_bh30_w103_3 & heap_bh30_w103_2;
      Compressor_bh30_176: Compressor_6_3
      port map ( R => CompressorOut_bh30_176_176,
                 X0 => CompressorIn_bh30_176_290);
   heap_bh30_w103_10 <= CompressorOut_bh30_176_176(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w104_9 <= CompressorOut_bh30_176_176(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w105_8 <= CompressorOut_bh30_176_176(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_177_291 <= heap_bh30_w104_7 & heap_bh30_w104_6 & heap_bh30_w104_5 & heap_bh30_w104_4 & heap_bh30_w104_3 & heap_bh30_w104_2;
      Compressor_bh30_177: Compressor_6_3
      port map ( R => CompressorOut_bh30_177_177,
                 X0 => CompressorIn_bh30_177_291);
   heap_bh30_w104_10 <= CompressorOut_bh30_177_177(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w105_9 <= CompressorOut_bh30_177_177(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w106_8 <= CompressorOut_bh30_177_177(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_178_292 <= heap_bh30_w105_7 & heap_bh30_w105_6 & heap_bh30_w105_5 & heap_bh30_w105_4 & heap_bh30_w105_3 & heap_bh30_w105_2;
      Compressor_bh30_178: Compressor_6_3
      port map ( R => CompressorOut_bh30_178_178,
                 X0 => CompressorIn_bh30_178_292);
   heap_bh30_w105_10 <= CompressorOut_bh30_178_178(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w106_9 <= CompressorOut_bh30_178_178(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w107_8 <= CompressorOut_bh30_178_178(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_179_293 <= heap_bh30_w106_7 & heap_bh30_w106_6 & heap_bh30_w106_5 & heap_bh30_w106_4 & heap_bh30_w106_3 & heap_bh30_w106_2;
      Compressor_bh30_179: Compressor_6_3
      port map ( R => CompressorOut_bh30_179_179,
                 X0 => CompressorIn_bh30_179_293);
   heap_bh30_w106_10 <= CompressorOut_bh30_179_179(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w107_9 <= CompressorOut_bh30_179_179(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w108_7 <= CompressorOut_bh30_179_179(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_180_294 <= heap_bh30_w107_7 & heap_bh30_w107_6 & heap_bh30_w107_5 & heap_bh30_w107_4 & heap_bh30_w107_3 & heap_bh30_w107_2;
      Compressor_bh30_180: Compressor_6_3
      port map ( R => CompressorOut_bh30_180_180,
                 X0 => CompressorIn_bh30_180_294);
   heap_bh30_w107_10 <= CompressorOut_bh30_180_180(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w108_8 <= CompressorOut_bh30_180_180(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w109_7 <= CompressorOut_bh30_180_180(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_181_295 <= heap_bh30_w108_6 & heap_bh30_w108_5 & heap_bh30_w108_4 & heap_bh30_w108_3 & heap_bh30_w108_2 & heap_bh30_w108_1;
      Compressor_bh30_181: Compressor_6_3
      port map ( R => CompressorOut_bh30_181_181,
                 X0 => CompressorIn_bh30_181_295);
   heap_bh30_w108_9 <= CompressorOut_bh30_181_181(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w109_8 <= CompressorOut_bh30_181_181(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w110_7 <= CompressorOut_bh30_181_181(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_182_296 <= heap_bh30_w109_6 & heap_bh30_w109_5 & heap_bh30_w109_4 & heap_bh30_w109_3 & heap_bh30_w109_2 & heap_bh30_w109_1;
      Compressor_bh30_182: Compressor_6_3
      port map ( R => CompressorOut_bh30_182_182,
                 X0 => CompressorIn_bh30_182_296);
   heap_bh30_w109_9 <= CompressorOut_bh30_182_182(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w110_8 <= CompressorOut_bh30_182_182(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w111_7 <= CompressorOut_bh30_182_182(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_183_297 <= heap_bh30_w110_6 & heap_bh30_w110_5 & heap_bh30_w110_4 & heap_bh30_w110_3 & heap_bh30_w110_2 & heap_bh30_w110_1;
      Compressor_bh30_183: Compressor_6_3
      port map ( R => CompressorOut_bh30_183_183,
                 X0 => CompressorIn_bh30_183_297);
   heap_bh30_w110_9 <= CompressorOut_bh30_183_183(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w111_8 <= CompressorOut_bh30_183_183(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w112_6 <= CompressorOut_bh30_183_183(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_184_298 <= heap_bh30_w111_6 & heap_bh30_w111_5 & heap_bh30_w111_4 & heap_bh30_w111_3 & heap_bh30_w111_2 & heap_bh30_w111_1;
      Compressor_bh30_184: Compressor_6_3
      port map ( R => CompressorOut_bh30_184_184,
                 X0 => CompressorIn_bh30_184_298);
   heap_bh30_w111_9 <= CompressorOut_bh30_184_184(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w112_7 <= CompressorOut_bh30_184_184(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w113_6 <= CompressorOut_bh30_184_184(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_185_299 <= heap_bh30_w112_5 & heap_bh30_w112_4 & heap_bh30_w112_3 & heap_bh30_w112_2 & heap_bh30_w112_1 & heap_bh30_w112_0;
      Compressor_bh30_185: Compressor_6_3
      port map ( R => CompressorOut_bh30_185_185,
                 X0 => CompressorIn_bh30_185_299);
   heap_bh30_w112_8 <= CompressorOut_bh30_185_185(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w113_7 <= CompressorOut_bh30_185_185(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w114_6 <= CompressorOut_bh30_185_185(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_186_300 <= heap_bh30_w113_5 & heap_bh30_w113_4 & heap_bh30_w113_3 & heap_bh30_w113_2 & heap_bh30_w113_1 & heap_bh30_w113_0;
      Compressor_bh30_186: Compressor_6_3
      port map ( R => CompressorOut_bh30_186_186,
                 X0 => CompressorIn_bh30_186_300);
   heap_bh30_w113_8 <= CompressorOut_bh30_186_186(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w114_7 <= CompressorOut_bh30_186_186(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w115_6 <= CompressorOut_bh30_186_186(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_187_301 <= heap_bh30_w114_5 & heap_bh30_w114_4 & heap_bh30_w114_3 & heap_bh30_w114_2 & heap_bh30_w114_1 & heap_bh30_w114_0;
      Compressor_bh30_187: Compressor_6_3
      port map ( R => CompressorOut_bh30_187_187,
                 X0 => CompressorIn_bh30_187_301);
   heap_bh30_w114_8 <= CompressorOut_bh30_187_187(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w115_7 <= CompressorOut_bh30_187_187(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w116_6 <= CompressorOut_bh30_187_187(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_188_302 <= heap_bh30_w115_5 & heap_bh30_w115_4 & heap_bh30_w115_3 & heap_bh30_w115_2 & heap_bh30_w115_1 & heap_bh30_w115_0;
      Compressor_bh30_188: Compressor_6_3
      port map ( R => CompressorOut_bh30_188_188,
                 X0 => CompressorIn_bh30_188_302);
   heap_bh30_w115_8 <= CompressorOut_bh30_188_188(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w116_7 <= CompressorOut_bh30_188_188(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w117_6 <= CompressorOut_bh30_188_188(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_189_303 <= heap_bh30_w116_5 & heap_bh30_w116_4 & heap_bh30_w116_3 & heap_bh30_w116_2 & heap_bh30_w116_1 & heap_bh30_w116_0;
      Compressor_bh30_189: Compressor_6_3
      port map ( R => CompressorOut_bh30_189_189,
                 X0 => CompressorIn_bh30_189_303);
   heap_bh30_w116_8 <= CompressorOut_bh30_189_189(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w117_7 <= CompressorOut_bh30_189_189(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w118_6 <= CompressorOut_bh30_189_189(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_190_304 <= heap_bh30_w117_5 & heap_bh30_w117_4 & heap_bh30_w117_3 & heap_bh30_w117_2 & heap_bh30_w117_1 & heap_bh30_w117_0;
      Compressor_bh30_190: Compressor_6_3
      port map ( R => CompressorOut_bh30_190_190,
                 X0 => CompressorIn_bh30_190_304);
   heap_bh30_w117_8 <= CompressorOut_bh30_190_190(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w118_7 <= CompressorOut_bh30_190_190(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w119_6 <= CompressorOut_bh30_190_190(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_191_305 <= heap_bh30_w118_5 & heap_bh30_w118_4 & heap_bh30_w118_3 & heap_bh30_w118_2 & heap_bh30_w118_1 & heap_bh30_w118_0;
      Compressor_bh30_191: Compressor_6_3
      port map ( R => CompressorOut_bh30_191_191,
                 X0 => CompressorIn_bh30_191_305);
   heap_bh30_w118_8 <= CompressorOut_bh30_191_191(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w119_7 <= CompressorOut_bh30_191_191(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w120_6 <= CompressorOut_bh30_191_191(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_192_306 <= heap_bh30_w119_5 & heap_bh30_w119_4 & heap_bh30_w119_3 & heap_bh30_w119_2 & heap_bh30_w119_1 & heap_bh30_w119_0;
      Compressor_bh30_192: Compressor_6_3
      port map ( R => CompressorOut_bh30_192_192,
                 X0 => CompressorIn_bh30_192_306);
   heap_bh30_w119_8 <= CompressorOut_bh30_192_192(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w120_7 <= CompressorOut_bh30_192_192(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w121_6 <= CompressorOut_bh30_192_192(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_193_307 <= heap_bh30_w120_5 & heap_bh30_w120_4 & heap_bh30_w120_3 & heap_bh30_w120_2 & heap_bh30_w120_1 & heap_bh30_w120_0;
      Compressor_bh30_193: Compressor_6_3
      port map ( R => CompressorOut_bh30_193_193,
                 X0 => CompressorIn_bh30_193_307);
   heap_bh30_w120_8 <= CompressorOut_bh30_193_193(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w121_7 <= CompressorOut_bh30_193_193(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w122_6 <= CompressorOut_bh30_193_193(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_194_308 <= heap_bh30_w121_5 & heap_bh30_w121_4 & heap_bh30_w121_3 & heap_bh30_w121_2 & heap_bh30_w121_1 & heap_bh30_w121_0;
      Compressor_bh30_194: Compressor_6_3
      port map ( R => CompressorOut_bh30_194_194,
                 X0 => CompressorIn_bh30_194_308);
   heap_bh30_w121_8 <= CompressorOut_bh30_194_194(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w122_7 <= CompressorOut_bh30_194_194(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w123_6 <= CompressorOut_bh30_194_194(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_195_309 <= heap_bh30_w122_5 & heap_bh30_w122_4 & heap_bh30_w122_3 & heap_bh30_w122_2 & heap_bh30_w122_1 & heap_bh30_w122_0;
      Compressor_bh30_195: Compressor_6_3
      port map ( R => CompressorOut_bh30_195_195,
                 X0 => CompressorIn_bh30_195_309);
   heap_bh30_w122_8 <= CompressorOut_bh30_195_195(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w123_7 <= CompressorOut_bh30_195_195(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w124_6 <= CompressorOut_bh30_195_195(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_196_310 <= heap_bh30_w123_5 & heap_bh30_w123_4 & heap_bh30_w123_3 & heap_bh30_w123_2 & heap_bh30_w123_1 & heap_bh30_w123_0;
      Compressor_bh30_196: Compressor_6_3
      port map ( R => CompressorOut_bh30_196_196,
                 X0 => CompressorIn_bh30_196_310);
   heap_bh30_w123_8 <= CompressorOut_bh30_196_196(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w124_7 <= CompressorOut_bh30_196_196(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w125_6 <= CompressorOut_bh30_196_196(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_197_311 <= heap_bh30_w124_5 & heap_bh30_w124_4 & heap_bh30_w124_3 & heap_bh30_w124_2 & heap_bh30_w124_1 & heap_bh30_w124_0;
      Compressor_bh30_197: Compressor_6_3
      port map ( R => CompressorOut_bh30_197_197,
                 X0 => CompressorIn_bh30_197_311);
   heap_bh30_w124_8 <= CompressorOut_bh30_197_197(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w125_7 <= CompressorOut_bh30_197_197(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w126_6 <= CompressorOut_bh30_197_197(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_198_312 <= heap_bh30_w125_5 & heap_bh30_w125_4 & heap_bh30_w125_3 & heap_bh30_w125_2 & heap_bh30_w125_1 & heap_bh30_w125_0;
      Compressor_bh30_198: Compressor_6_3
      port map ( R => CompressorOut_bh30_198_198,
                 X0 => CompressorIn_bh30_198_312);
   heap_bh30_w125_8 <= CompressorOut_bh30_198_198(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w126_7 <= CompressorOut_bh30_198_198(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w127_6 <= CompressorOut_bh30_198_198(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_199_313 <= heap_bh30_w126_5 & heap_bh30_w126_4 & heap_bh30_w126_3 & heap_bh30_w126_2 & heap_bh30_w126_1 & heap_bh30_w126_0;
      Compressor_bh30_199: Compressor_6_3
      port map ( R => CompressorOut_bh30_199_199,
                 X0 => CompressorIn_bh30_199_313);
   heap_bh30_w126_8 <= CompressorOut_bh30_199_199(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w127_7 <= CompressorOut_bh30_199_199(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w128_6 <= CompressorOut_bh30_199_199(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_200_314 <= heap_bh30_w127_5 & heap_bh30_w127_4 & heap_bh30_w127_3 & heap_bh30_w127_2 & heap_bh30_w127_1 & heap_bh30_w127_0;
      Compressor_bh30_200: Compressor_6_3
      port map ( R => CompressorOut_bh30_200_200,
                 X0 => CompressorIn_bh30_200_314);
   heap_bh30_w127_8 <= CompressorOut_bh30_200_200(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w128_7 <= CompressorOut_bh30_200_200(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w129_5 <= CompressorOut_bh30_200_200(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_201_315 <= heap_bh30_w128_5 & heap_bh30_w128_4 & heap_bh30_w128_3 & heap_bh30_w128_2 & heap_bh30_w128_1 & heap_bh30_w128_0;
      Compressor_bh30_201: Compressor_6_3
      port map ( R => CompressorOut_bh30_201_201,
                 X0 => CompressorIn_bh30_201_315);
   heap_bh30_w128_8 <= CompressorOut_bh30_201_201(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w129_6 <= CompressorOut_bh30_201_201(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w130_5 <= CompressorOut_bh30_201_201(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_202_316 <= heap_bh30_w18_8 & heap_bh30_w18_9 & heap_bh30_w18_5 & heap_bh30_w18_4;
   CompressorIn_bh30_202_317(0) <= heap_bh30_w19_9;
      Compressor_bh30_202: Compressor_14_3
      port map ( R => CompressorOut_bh30_202_202,
                 X0 => CompressorIn_bh30_202_316,
                 X1 => CompressorIn_bh30_202_317);
   heap_bh30_w18_10 <= CompressorOut_bh30_202_202(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w19_10 <= CompressorOut_bh30_202_202(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w20_9 <= CompressorOut_bh30_202_202(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_203_318 <= heap_bh30_w21_8 & heap_bh30_w21_9 & heap_bh30_w21_5 & heap_bh30_w21_4;
   CompressorIn_bh30_203_319(0) <= heap_bh30_w22_9;
      Compressor_bh30_203: Compressor_14_3
      port map ( R => CompressorOut_bh30_203_203,
                 X0 => CompressorIn_bh30_203_318,
                 X1 => CompressorIn_bh30_203_319);
   heap_bh30_w21_10 <= CompressorOut_bh30_203_203(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w22_10 <= CompressorOut_bh30_203_203(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w23_10 <= CompressorOut_bh30_203_203(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_204_320 <= heap_bh30_w23_9 & heap_bh30_w23_5 & heap_bh30_w23_4 & heap_bh30_w23_3;
   CompressorIn_bh30_204_321(0) <= heap_bh30_w24_9;
      Compressor_bh30_204: Compressor_14_3
      port map ( R => CompressorOut_bh30_204_204,
                 X0 => CompressorIn_bh30_204_320,
                 X1 => CompressorIn_bh30_204_321);
   heap_bh30_w23_11 <= CompressorOut_bh30_204_204(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w24_11 <= CompressorOut_bh30_204_204(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w25_11 <= CompressorOut_bh30_204_204(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_205_322 <= heap_bh30_w24_10 & heap_bh30_w24_6 & heap_bh30_w24_5 & heap_bh30_w24_4;
   CompressorIn_bh30_205_323(0) <= heap_bh30_w25_10;
      Compressor_bh30_205: Compressor_14_3
      port map ( R => CompressorOut_bh30_205_205,
                 X0 => CompressorIn_bh30_205_322,
                 X1 => CompressorIn_bh30_205_323);
   heap_bh30_w24_12 <= CompressorOut_bh30_205_205(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w25_12 <= CompressorOut_bh30_205_205(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w26_10 <= CompressorOut_bh30_205_205(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_206_324 <= heap_bh30_w26_9 & heap_bh30_w26_5 & heap_bh30_w26_4 & heap_bh30_w26_3;
   CompressorIn_bh30_206_325(0) <= heap_bh30_w27_9;
      Compressor_bh30_206: Compressor_14_3
      port map ( R => CompressorOut_bh30_206_206,
                 X0 => CompressorIn_bh30_206_324,
                 X1 => CompressorIn_bh30_206_325);
   heap_bh30_w26_11 <= CompressorOut_bh30_206_206(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w27_11 <= CompressorOut_bh30_206_206(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w28_11 <= CompressorOut_bh30_206_206(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_207_326 <= heap_bh30_w27_10 & heap_bh30_w27_6 & heap_bh30_w27_5 & heap_bh30_w27_4;
   CompressorIn_bh30_207_327(0) <= heap_bh30_w28_10;
      Compressor_bh30_207: Compressor_14_3
      port map ( R => CompressorOut_bh30_207_207,
                 X0 => CompressorIn_bh30_207_326,
                 X1 => CompressorIn_bh30_207_327);
   heap_bh30_w27_12 <= CompressorOut_bh30_207_207(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w28_12 <= CompressorOut_bh30_207_207(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w29_10 <= CompressorOut_bh30_207_207(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_208_328 <= heap_bh30_w29_9 & heap_bh30_w29_5 & heap_bh30_w29_4 & heap_bh30_w29_3;
   CompressorIn_bh30_208_329(0) <= heap_bh30_w30_9;
      Compressor_bh30_208: Compressor_14_3
      port map ( R => CompressorOut_bh30_208_208,
                 X0 => CompressorIn_bh30_208_328,
                 X1 => CompressorIn_bh30_208_329);
   heap_bh30_w29_11 <= CompressorOut_bh30_208_208(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w30_11 <= CompressorOut_bh30_208_208(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w31_11 <= CompressorOut_bh30_208_208(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_209_330 <= heap_bh30_w30_10 & heap_bh30_w30_6 & heap_bh30_w30_5 & heap_bh30_w30_4;
   CompressorIn_bh30_209_331(0) <= heap_bh30_w31_10;
      Compressor_bh30_209: Compressor_14_3
      port map ( R => CompressorOut_bh30_209_209,
                 X0 => CompressorIn_bh30_209_330,
                 X1 => CompressorIn_bh30_209_331);
   heap_bh30_w30_12 <= CompressorOut_bh30_209_209(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w31_12 <= CompressorOut_bh30_209_209(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w32_10 <= CompressorOut_bh30_209_209(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_210_332 <= heap_bh30_w34_11 & heap_bh30_w34_7 & heap_bh30_w34_6 & heap_bh30_w34_5;
   CompressorIn_bh30_210_333(0) <= heap_bh30_w35_10;
      Compressor_bh30_210: Compressor_14_3
      port map ( R => CompressorOut_bh30_210_210,
                 X0 => CompressorIn_bh30_210_332,
                 X1 => CompressorIn_bh30_210_333);
   heap_bh30_w34_13 <= CompressorOut_bh30_210_210(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w35_12 <= CompressorOut_bh30_210_210(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w36_13 <= CompressorOut_bh30_210_210(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_211_334 <= heap_bh30_w37_11 & heap_bh30_w37_7 & heap_bh30_w37_6 & heap_bh30_w37_5;
   CompressorIn_bh30_211_335(0) <= heap_bh30_w38_10;
      Compressor_bh30_211: Compressor_14_3
      port map ( R => CompressorOut_bh30_211_211,
                 X0 => CompressorIn_bh30_211_334,
                 X1 => CompressorIn_bh30_211_335);
   heap_bh30_w37_13 <= CompressorOut_bh30_211_211(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w38_12 <= CompressorOut_bh30_211_211(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w39_13 <= CompressorOut_bh30_211_211(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_212_336 <= heap_bh30_w40_11 & heap_bh30_w40_7 & heap_bh30_w40_6 & heap_bh30_w40_5;
   CompressorIn_bh30_212_337(0) <= heap_bh30_w41_10;
      Compressor_bh30_212: Compressor_14_3
      port map ( R => CompressorOut_bh30_212_212,
                 X0 => CompressorIn_bh30_212_336,
                 X1 => CompressorIn_bh30_212_337);
   heap_bh30_w40_13 <= CompressorOut_bh30_212_212(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w41_12 <= CompressorOut_bh30_212_212(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w42_13 <= CompressorOut_bh30_212_212(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_213_338 <= heap_bh30_w43_11 & heap_bh30_w43_7 & heap_bh30_w43_6 & heap_bh30_w43_5;
   CompressorIn_bh30_213_339(0) <= heap_bh30_w44_10;
      Compressor_bh30_213: Compressor_14_3
      port map ( R => CompressorOut_bh30_213_213,
                 X0 => CompressorIn_bh30_213_338,
                 X1 => CompressorIn_bh30_213_339);
   heap_bh30_w43_13 <= CompressorOut_bh30_213_213(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w44_12 <= CompressorOut_bh30_213_213(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w45_13 <= CompressorOut_bh30_213_213(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_214_340 <= heap_bh30_w72_7 & heap_bh30_w72_6 & heap_bh30_w72_5 & heap_bh30_w72_4;
   CompressorIn_bh30_214_341(0) <= heap_bh30_w73_6;
      Compressor_bh30_214: Compressor_14_3
      port map ( R => CompressorOut_bh30_214_214,
                 X0 => CompressorIn_bh30_214_340,
                 X1 => CompressorIn_bh30_214_341);
   heap_bh30_w72_19 <= CompressorOut_bh30_214_214(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w73_19 <= CompressorOut_bh30_214_214(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w74_18 <= CompressorOut_bh30_214_214(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_215_342 <= heap_bh30_w75_7 & heap_bh30_w75_6 & heap_bh30_w75_5 & heap_bh30_w75_4;
   CompressorIn_bh30_215_343(0) <= heap_bh30_w76_6;
      Compressor_bh30_215: Compressor_14_3
      port map ( R => CompressorOut_bh30_215_215,
                 X0 => CompressorIn_bh30_215_342,
                 X1 => CompressorIn_bh30_215_343);
   heap_bh30_w75_19 <= CompressorOut_bh30_215_215(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w76_19 <= CompressorOut_bh30_215_215(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w77_18 <= CompressorOut_bh30_215_215(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_216_344 <= heap_bh30_w78_7 & heap_bh30_w78_6 & heap_bh30_w78_5 & heap_bh30_w78_4;
   CompressorIn_bh30_216_345(0) <= heap_bh30_w79_6;
      Compressor_bh30_216: Compressor_14_3
      port map ( R => CompressorOut_bh30_216_216,
                 X0 => CompressorIn_bh30_216_344,
                 X1 => CompressorIn_bh30_216_345);
   heap_bh30_w78_19 <= CompressorOut_bh30_216_216(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w79_19 <= CompressorOut_bh30_216_216(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w80_18 <= CompressorOut_bh30_216_216(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_217_346 <= heap_bh30_w81_7 & heap_bh30_w81_6 & heap_bh30_w81_5 & heap_bh30_w81_4;
   CompressorIn_bh30_217_347(0) <= heap_bh30_w82_6;
      Compressor_bh30_217: Compressor_14_3
      port map ( R => CompressorOut_bh30_217_217,
                 X0 => CompressorIn_bh30_217_346,
                 X1 => CompressorIn_bh30_217_347);
   heap_bh30_w81_19 <= CompressorOut_bh30_217_217(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w82_19 <= CompressorOut_bh30_217_217(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w83_18 <= CompressorOut_bh30_217_217(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_218_348 <= heap_bh30_w84_7 & heap_bh30_w84_6 & heap_bh30_w84_5 & heap_bh30_w84_4;
   CompressorIn_bh30_218_349(0) <= heap_bh30_w85_6;
      Compressor_bh30_218: Compressor_14_3
      port map ( R => CompressorOut_bh30_218_218,
                 X0 => CompressorIn_bh30_218_348,
                 X1 => CompressorIn_bh30_218_349);
   heap_bh30_w84_19 <= CompressorOut_bh30_218_218(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w85_19 <= CompressorOut_bh30_218_218(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w86_18 <= CompressorOut_bh30_218_218(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_219_350 <= heap_bh30_w87_7 & heap_bh30_w87_6 & heap_bh30_w87_5 & heap_bh30_w87_4;
   CompressorIn_bh30_219_351(0) <= heap_bh30_w88_6;
      Compressor_bh30_219: Compressor_14_3
      port map ( R => CompressorOut_bh30_219_219,
                 X0 => CompressorIn_bh30_219_350,
                 X1 => CompressorIn_bh30_219_351);
   heap_bh30_w87_19 <= CompressorOut_bh30_219_219(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w88_19 <= CompressorOut_bh30_219_219(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w89_18 <= CompressorOut_bh30_219_219(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_220_352 <= heap_bh30_w90_6 & heap_bh30_w90_5 & heap_bh30_w90_4 & heap_bh30_w90_3;
   CompressorIn_bh30_220_353(0) <= heap_bh30_w91_5;
      Compressor_bh30_220: Compressor_14_3
      port map ( R => CompressorOut_bh30_220_220,
                 X0 => CompressorIn_bh30_220_352,
                 X1 => CompressorIn_bh30_220_353);
   heap_bh30_w90_18 <= CompressorOut_bh30_220_220(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w91_17 <= CompressorOut_bh30_220_220(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w92_14 <= CompressorOut_bh30_220_220(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_221_354 <= heap_bh30_w93_4 & heap_bh30_w93_3 & heap_bh30_w93_2 & heap_bh30_w93_1;
   CompressorIn_bh30_221_355(0) <= heap_bh30_w94_3;
      Compressor_bh30_221: Compressor_14_3
      port map ( R => CompressorOut_bh30_221_221,
                 X0 => CompressorIn_bh30_221_354,
                 X1 => CompressorIn_bh30_221_355);
   heap_bh30_w93_13 <= CompressorOut_bh30_221_221(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w94_12 <= CompressorOut_bh30_221_221(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w95_11 <= CompressorOut_bh30_221_221(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_222_356 <= heap_bh30_w129_4 & heap_bh30_w129_3 & heap_bh30_w129_2 & heap_bh30_w129_1;
   CompressorIn_bh30_222_357(0) <= heap_bh30_w130_4;
      Compressor_bh30_222: Compressor_14_3
      port map ( R => CompressorOut_bh30_222_222,
                 X0 => CompressorIn_bh30_222_356,
                 X1 => CompressorIn_bh30_222_357);
   heap_bh30_w129_7 <= CompressorOut_bh30_222_222(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w130_6 <= CompressorOut_bh30_222_222(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w131_5 <= CompressorOut_bh30_222_222(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_223_358 <= heap_bh30_w130_3 & heap_bh30_w130_2 & heap_bh30_w130_1 & heap_bh30_w130_0;
   CompressorIn_bh30_223_359(0) <= heap_bh30_w131_4;
      Compressor_bh30_223: Compressor_14_3
      port map ( R => CompressorOut_bh30_223_223,
                 X0 => CompressorIn_bh30_223_358,
                 X1 => CompressorIn_bh30_223_359);
   heap_bh30_w130_7 <= CompressorOut_bh30_223_223(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w131_6 <= CompressorOut_bh30_223_223(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w132_4 <= CompressorOut_bh30_223_223(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_224_360 <= heap_bh30_w131_3 & heap_bh30_w131_2 & heap_bh30_w131_1 & heap_bh30_w131_0;
   CompressorIn_bh30_224_361(0) <= heap_bh30_w132_3;
      Compressor_bh30_224: Compressor_14_3
      port map ( R => CompressorOut_bh30_224_224,
                 X0 => CompressorIn_bh30_224_360,
                 X1 => CompressorIn_bh30_224_361);
   heap_bh30_w131_7 <= CompressorOut_bh30_224_224(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w132_5 <= CompressorOut_bh30_224_224(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w133_4 <= CompressorOut_bh30_224_224(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_225_362 <= heap_bh30_w133_3 & heap_bh30_w133_2 & heap_bh30_w133_1 & heap_bh30_w133_0;
   CompressorIn_bh30_225_363(0) <= heap_bh30_w134_3;
      Compressor_bh30_225: Compressor_14_3
      port map ( R => CompressorOut_bh30_225_225,
                 X0 => CompressorIn_bh30_225_362,
                 X1 => CompressorIn_bh30_225_363);
   heap_bh30_w133_5 <= CompressorOut_bh30_225_225(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w134_4 <= CompressorOut_bh30_225_225(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w135_4 <= CompressorOut_bh30_225_225(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_226_364 <= heap_bh30_w135_3 & heap_bh30_w135_2 & heap_bh30_w135_1 & heap_bh30_w135_0;
   CompressorIn_bh30_226_365(0) <= heap_bh30_w136_3;
      Compressor_bh30_226: Compressor_14_3
      port map ( R => CompressorOut_bh30_226_226,
                 X0 => CompressorIn_bh30_226_364,
                 X1 => CompressorIn_bh30_226_365);
   heap_bh30_w135_5 <= CompressorOut_bh30_226_226(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w136_4 <= CompressorOut_bh30_226_226(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w137_4 <= CompressorOut_bh30_226_226(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_227_366 <= heap_bh30_w137_3 & heap_bh30_w137_2 & heap_bh30_w137_1 & heap_bh30_w137_0;
   CompressorIn_bh30_227_367(0) <= heap_bh30_w138_3;
      Compressor_bh30_227: Compressor_14_3
      port map ( R => CompressorOut_bh30_227_227,
                 X0 => CompressorIn_bh30_227_366,
                 X1 => CompressorIn_bh30_227_367);
   heap_bh30_w137_5 <= CompressorOut_bh30_227_227(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w138_4 <= CompressorOut_bh30_227_227(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w139_4 <= CompressorOut_bh30_227_227(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_228_368 <= heap_bh30_w139_3 & heap_bh30_w139_2 & heap_bh30_w139_1 & heap_bh30_w139_0;
   CompressorIn_bh30_228_369(0) <= heap_bh30_w140_3;
      Compressor_bh30_228: Compressor_14_3
      port map ( R => CompressorOut_bh30_228_228,
                 X0 => CompressorIn_bh30_228_368,
                 X1 => CompressorIn_bh30_228_369);
   heap_bh30_w139_5 <= CompressorOut_bh30_228_228(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w140_4 <= CompressorOut_bh30_228_228(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w141_4 <= CompressorOut_bh30_228_228(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_229_370 <= heap_bh30_w141_3 & heap_bh30_w141_2 & heap_bh30_w141_1 & heap_bh30_w141_0;
   CompressorIn_bh30_229_371(0) <= heap_bh30_w142_3;
      Compressor_bh30_229: Compressor_14_3
      port map ( R => CompressorOut_bh30_229_229,
                 X0 => CompressorIn_bh30_229_370,
                 X1 => CompressorIn_bh30_229_371);
   heap_bh30_w141_5 <= CompressorOut_bh30_229_229(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w142_4 <= CompressorOut_bh30_229_229(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w143_4 <= CompressorOut_bh30_229_229(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_230_372 <= heap_bh30_w143_3 & heap_bh30_w143_2 & heap_bh30_w143_1 & heap_bh30_w143_0;
   CompressorIn_bh30_230_373(0) <= heap_bh30_w144_3;
      Compressor_bh30_230: Compressor_14_3
      port map ( R => CompressorOut_bh30_230_230,
                 X0 => CompressorIn_bh30_230_372,
                 X1 => CompressorIn_bh30_230_373);
   heap_bh30_w143_5 <= CompressorOut_bh30_230_230(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w144_4 <= CompressorOut_bh30_230_230(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w145_4 <= CompressorOut_bh30_230_230(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_231_374 <= heap_bh30_w145_3 & heap_bh30_w145_2 & heap_bh30_w145_1 & heap_bh30_w145_0;
   CompressorIn_bh30_231_375(0) <= heap_bh30_w146_2;
      Compressor_bh30_231: Compressor_14_3
      port map ( R => CompressorOut_bh30_231_231,
                 X0 => CompressorIn_bh30_231_374,
                 X1 => CompressorIn_bh30_231_375);
   heap_bh30_w145_5 <= CompressorOut_bh30_231_231(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w146_3 <= CompressorOut_bh30_231_231(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w147_3 <= CompressorOut_bh30_231_231(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_232_376 <= heap_bh30_w46_11 & heap_bh30_w46_7 & heap_bh30_w46_6 & heap_bh30_w46_5 & heap_bh30_w46_4;
      Compressor_bh30_232: Compressor_5_3
      port map ( R => CompressorOut_bh30_232_232,
                 X0 => CompressorIn_bh30_232_376);
   heap_bh30_w46_13 <= CompressorOut_bh30_232_232(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w47_14 <= CompressorOut_bh30_232_232(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w48_15 <= CompressorOut_bh30_232_232(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_233_377 <= heap_bh30_w32_9 & heap_bh30_w32_5 & heap_bh30_w32_4 & heap_bh30_w32_3;
      Compressor_bh30_233: Compressor_4_3
      port map ( R => CompressorOut_bh30_233_233,
                 X0 => CompressorIn_bh30_233_377);
   heap_bh30_w32_11 <= CompressorOut_bh30_233_233(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w33_13 <= CompressorOut_bh30_233_233(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w34_14 <= CompressorOut_bh30_233_233(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_234_378 <= heap_bh30_w35_6 & heap_bh30_w35_5 & heap_bh30_w35_4 & heap_bh30_w35_3;
      Compressor_bh30_234: Compressor_4_3
      port map ( R => CompressorOut_bh30_234_234,
                 X0 => CompressorIn_bh30_234_378);
   heap_bh30_w35_13 <= CompressorOut_bh30_234_234(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w36_14 <= CompressorOut_bh30_234_234(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w37_14 <= CompressorOut_bh30_234_234(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_235_379 <= heap_bh30_w38_6 & heap_bh30_w38_5 & heap_bh30_w38_4 & heap_bh30_w38_3;
      Compressor_bh30_235: Compressor_4_3
      port map ( R => CompressorOut_bh30_235_235,
                 X0 => CompressorIn_bh30_235_379);
   heap_bh30_w38_13 <= CompressorOut_bh30_235_235(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w39_14 <= CompressorOut_bh30_235_235(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w40_14 <= CompressorOut_bh30_235_235(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_236_380 <= heap_bh30_w41_6 & heap_bh30_w41_5 & heap_bh30_w41_4 & heap_bh30_w41_3;
      Compressor_bh30_236: Compressor_4_3
      port map ( R => CompressorOut_bh30_236_236,
                 X0 => CompressorIn_bh30_236_380);
   heap_bh30_w41_13 <= CompressorOut_bh30_236_236(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w42_14 <= CompressorOut_bh30_236_236(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w43_14 <= CompressorOut_bh30_236_236(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_237_381 <= heap_bh30_w44_6 & heap_bh30_w44_5 & heap_bh30_w44_4 & heap_bh30_w44_3;
      Compressor_bh30_237: Compressor_4_3
      port map ( R => CompressorOut_bh30_237_237,
                 X0 => CompressorIn_bh30_237_381);
   heap_bh30_w44_13 <= CompressorOut_bh30_237_237(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w45_14 <= CompressorOut_bh30_237_237(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w46_14 <= CompressorOut_bh30_237_237(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_238_382 <= heap_bh30_w2_1 & heap_bh30_w2_0 & heap_bh30_w2_2;
   CompressorIn_bh30_238_383 <= heap_bh30_w3_4 & heap_bh30_w3_3;
      Compressor_bh30_238: Compressor_23_3
      port map ( R => CompressorOut_bh30_238_238,
                 X0 => CompressorIn_bh30_238_382,
                 X1 => CompressorIn_bh30_238_383);
   heap_bh30_w2_3 <= CompressorOut_bh30_238_238(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w3_5 <= CompressorOut_bh30_238_238(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w4_5 <= CompressorOut_bh30_238_238(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_239_384 <= heap_bh30_w4_0 & heap_bh30_w4_4 & heap_bh30_w4_3;
   CompressorIn_bh30_239_385 <= heap_bh30_w5_5 & heap_bh30_w5_4;
      Compressor_bh30_239: Compressor_23_3
      port map ( R => CompressorOut_bh30_239_239,
                 X0 => CompressorIn_bh30_239_384,
                 X1 => CompressorIn_bh30_239_385);
   heap_bh30_w4_6 <= CompressorOut_bh30_239_239(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w5_6 <= CompressorOut_bh30_239_239(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w6_7 <= CompressorOut_bh30_239_239(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_240_386 <= heap_bh30_w6_6 & heap_bh30_w6_5 & heap_bh30_w6_4;
   CompressorIn_bh30_240_387 <= heap_bh30_w7_6 & heap_bh30_w7_5;
      Compressor_bh30_240: Compressor_23_3
      port map ( R => CompressorOut_bh30_240_240,
                 X0 => CompressorIn_bh30_240_386,
                 X1 => CompressorIn_bh30_240_387);
   heap_bh30_w6_8 <= CompressorOut_bh30_240_240(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w7_7 <= CompressorOut_bh30_240_240(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w8_7 <= CompressorOut_bh30_240_240(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_241_388 <= heap_bh30_w12_7 & heap_bh30_w12_8 & heap_bh30_w12_4;
   CompressorIn_bh30_241_389 <= heap_bh30_w13_8 & heap_bh30_w13_4;
      Compressor_bh30_241: Compressor_23_3
      port map ( R => CompressorOut_bh30_241_241,
                 X0 => CompressorIn_bh30_241_388,
                 X1 => CompressorIn_bh30_241_389);
   heap_bh30_w12_9 <= CompressorOut_bh30_241_241(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w13_9 <= CompressorOut_bh30_241_241(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w14_8 <= CompressorOut_bh30_241_241(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_242_390 <= heap_bh30_w15_7 & heap_bh30_w15_8 & heap_bh30_w15_4;
   CompressorIn_bh30_242_391 <= heap_bh30_w16_9 & heap_bh30_w16_5;
      Compressor_bh30_242: Compressor_23_3
      port map ( R => CompressorOut_bh30_242_242,
                 X0 => CompressorIn_bh30_242_390,
                 X1 => CompressorIn_bh30_242_391);
   heap_bh30_w15_9 <= CompressorOut_bh30_242_242(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w16_10 <= CompressorOut_bh30_242_242(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w17_9 <= CompressorOut_bh30_242_242(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_243_392 <= heap_bh30_w69_6 & heap_bh30_w69_5 & heap_bh30_w69_4;
   CompressorIn_bh30_243_393 <= heap_bh30_w70_5 & heap_bh30_w70_4;
      Compressor_bh30_243: Compressor_23_3
      port map ( R => CompressorOut_bh30_243_243,
                 X0 => CompressorIn_bh30_243_392,
                 X1 => CompressorIn_bh30_243_393);
   heap_bh30_w69_18 <= CompressorOut_bh30_243_243(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w70_18 <= CompressorOut_bh30_243_243(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w71_18 <= CompressorOut_bh30_243_243(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_244_394 <= heap_bh30_w147_2 & heap_bh30_w147_1 & heap_bh30_w147_0;
   CompressorIn_bh30_244_395 <= heap_bh30_w148_2 & heap_bh30_w148_1;
      Compressor_bh30_244: Compressor_23_3
      port map ( R => CompressorOut_bh30_244_244,
                 X0 => CompressorIn_bh30_244_394,
                 X1 => CompressorIn_bh30_244_395);
   heap_bh30_w147_4 <= CompressorOut_bh30_244_244(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w148_3 <= CompressorOut_bh30_244_244(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w149_3 <= CompressorOut_bh30_244_244(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_245_396 <= heap_bh30_w149_2 & heap_bh30_w149_1 & heap_bh30_w149_0;
   CompressorIn_bh30_245_397 <= heap_bh30_w150_2 & heap_bh30_w150_1;
      Compressor_bh30_245: Compressor_23_3
      port map ( R => CompressorOut_bh30_245_245,
                 X0 => CompressorIn_bh30_245_396,
                 X1 => CompressorIn_bh30_245_397);
   heap_bh30_w149_4 <= CompressorOut_bh30_245_245(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w150_3 <= CompressorOut_bh30_245_245(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w151_3 <= CompressorOut_bh30_245_245(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_246_398 <= heap_bh30_w151_2 & heap_bh30_w151_1 & heap_bh30_w151_0;
   CompressorIn_bh30_246_399 <= heap_bh30_w152_2 & heap_bh30_w152_1;
      Compressor_bh30_246: Compressor_23_3
      port map ( R => CompressorOut_bh30_246_246,
                 X0 => CompressorIn_bh30_246_398,
                 X1 => CompressorIn_bh30_246_399);
   heap_bh30_w151_4 <= CompressorOut_bh30_246_246(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w152_3 <= CompressorOut_bh30_246_246(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w153_3 <= CompressorOut_bh30_246_246(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_247_400 <= heap_bh30_w153_2 & heap_bh30_w153_1 & heap_bh30_w153_0;
   CompressorIn_bh30_247_401 <= heap_bh30_w154_2 & heap_bh30_w154_1;
      Compressor_bh30_247: Compressor_23_3
      port map ( R => CompressorOut_bh30_247_247,
                 X0 => CompressorIn_bh30_247_400,
                 X1 => CompressorIn_bh30_247_401);
   heap_bh30_w153_4 <= CompressorOut_bh30_247_247(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w154_3 <= CompressorOut_bh30_247_247(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w155_3 <= CompressorOut_bh30_247_247(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_248_402 <= heap_bh30_w155_2 & heap_bh30_w155_1 & heap_bh30_w155_0;
   CompressorIn_bh30_248_403 <= heap_bh30_w156_1 & heap_bh30_w156_0;
      Compressor_bh30_248: Compressor_23_3
      port map ( R => CompressorOut_bh30_248_248,
                 X0 => CompressorIn_bh30_248_402,
                 X1 => CompressorIn_bh30_248_403);
   heap_bh30_w155_4 <= CompressorOut_bh30_248_248(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w156_2 <= CompressorOut_bh30_248_248(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w157_2 <= CompressorOut_bh30_248_248(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_249_404 <= heap_bh30_w17_8 & heap_bh30_w17_4 & heap_bh30_w17_3;
      Compressor_bh30_249: Compressor_3_2
      port map ( R => CompressorOut_bh30_249_249,
                 X0 => CompressorIn_bh30_249_404);
   heap_bh30_w17_10 <= CompressorOut_bh30_249_249(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w18_11 <= CompressorOut_bh30_249_249(1); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_250_405 <= heap_bh30_w20_8 & heap_bh30_w20_4 & heap_bh30_w20_3;
      Compressor_bh30_250: Compressor_3_2
      port map ( R => CompressorOut_bh30_250_250,
                 X0 => CompressorIn_bh30_250_405);
   heap_bh30_w20_10 <= CompressorOut_bh30_250_250(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w21_11 <= CompressorOut_bh30_250_250(1); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_251_406 <= heap_bh30_w25_6 & heap_bh30_w25_5 & heap_bh30_w25_4;
      Compressor_bh30_251: Compressor_3_2
      port map ( R => CompressorOut_bh30_251_251,
                 X0 => CompressorIn_bh30_251_406);
   heap_bh30_w25_13 <= CompressorOut_bh30_251_251(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w26_12 <= CompressorOut_bh30_251_251(1); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_252_407 <= heap_bh30_w28_6 & heap_bh30_w28_5 & heap_bh30_w28_4;
      Compressor_bh30_252: Compressor_3_2
      port map ( R => CompressorOut_bh30_252_252,
                 X0 => CompressorIn_bh30_252_407);
   heap_bh30_w28_13 <= CompressorOut_bh30_252_252(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w29_12 <= CompressorOut_bh30_252_252(1); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_253_408 <= heap_bh30_w31_6 & heap_bh30_w31_5 & heap_bh30_w31_4;
      Compressor_bh30_253: Compressor_3_2
      port map ( R => CompressorOut_bh30_253_253,
                 X0 => CompressorIn_bh30_253_408);
   heap_bh30_w31_13 <= CompressorOut_bh30_253_253(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w32_12 <= CompressorOut_bh30_253_253(1); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_254_409 <= heap_bh30_w71_5 & heap_bh30_w71_4 & heap_bh30_w71_3;
      Compressor_bh30_254: Compressor_3_2
      port map ( R => CompressorOut_bh30_254_254,
                 X0 => CompressorIn_bh30_254_409);
   heap_bh30_w71_19 <= CompressorOut_bh30_254_254(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w72_20 <= CompressorOut_bh30_254_254(1); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_255_410 <= heap_bh30_w74_5 & heap_bh30_w74_4 & heap_bh30_w74_3;
      Compressor_bh30_255: Compressor_3_2
      port map ( R => CompressorOut_bh30_255_255,
                 X0 => CompressorIn_bh30_255_410);
   heap_bh30_w74_19 <= CompressorOut_bh30_255_255(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w75_20 <= CompressorOut_bh30_255_255(1); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_256_411 <= heap_bh30_w77_5 & heap_bh30_w77_4 & heap_bh30_w77_3;
      Compressor_bh30_256: Compressor_3_2
      port map ( R => CompressorOut_bh30_256_256,
                 X0 => CompressorIn_bh30_256_411);
   heap_bh30_w77_19 <= CompressorOut_bh30_256_256(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w78_20 <= CompressorOut_bh30_256_256(1); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_257_412 <= heap_bh30_w80_5 & heap_bh30_w80_4 & heap_bh30_w80_3;
      Compressor_bh30_257: Compressor_3_2
      port map ( R => CompressorOut_bh30_257_257,
                 X0 => CompressorIn_bh30_257_412);
   heap_bh30_w80_19 <= CompressorOut_bh30_257_257(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w81_20 <= CompressorOut_bh30_257_257(1); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_258_413 <= heap_bh30_w83_5 & heap_bh30_w83_4 & heap_bh30_w83_3;
      Compressor_bh30_258: Compressor_3_2
      port map ( R => CompressorOut_bh30_258_258,
                 X0 => CompressorIn_bh30_258_413);
   heap_bh30_w83_19 <= CompressorOut_bh30_258_258(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w84_20 <= CompressorOut_bh30_258_258(1); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_259_414 <= heap_bh30_w86_5 & heap_bh30_w86_4 & heap_bh30_w86_3;
      Compressor_bh30_259: Compressor_3_2
      port map ( R => CompressorOut_bh30_259_259,
                 X0 => CompressorIn_bh30_259_414);
   heap_bh30_w86_19 <= CompressorOut_bh30_259_259(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w87_20 <= CompressorOut_bh30_259_259(1); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_260_415 <= heap_bh30_w89_5 & heap_bh30_w89_4 & heap_bh30_w89_3;
      Compressor_bh30_260: Compressor_3_2
      port map ( R => CompressorOut_bh30_260_260,
                 X0 => CompressorIn_bh30_260_415);
   heap_bh30_w89_19 <= CompressorOut_bh30_260_260(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w90_19 <= CompressorOut_bh30_260_260(1); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_261_416 <= heap_bh30_w92_3 & heap_bh30_w92_2 & heap_bh30_w92_1;
      Compressor_bh30_261: Compressor_3_2
      port map ( R => CompressorOut_bh30_261_261,
                 X0 => CompressorIn_bh30_261_416);
   heap_bh30_w92_15 <= CompressorOut_bh30_261_261(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w93_14 <= CompressorOut_bh30_261_261(1); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_262_417 <= heap_bh30_w132_2 & heap_bh30_w132_1 & heap_bh30_w132_0;
      Compressor_bh30_262: Compressor_3_2
      port map ( R => CompressorOut_bh30_262_262,
                 X0 => CompressorIn_bh30_262_417);
   heap_bh30_w132_6 <= CompressorOut_bh30_262_262(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w133_6 <= CompressorOut_bh30_262_262(1); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_263_418 <= heap_bh30_w134_2 & heap_bh30_w134_1 & heap_bh30_w134_0;
      Compressor_bh30_263: Compressor_3_2
      port map ( R => CompressorOut_bh30_263_263,
                 X0 => CompressorIn_bh30_263_418);
   heap_bh30_w134_5 <= CompressorOut_bh30_263_263(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w135_6 <= CompressorOut_bh30_263_263(1); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_264_419 <= heap_bh30_w136_2 & heap_bh30_w136_1 & heap_bh30_w136_0;
      Compressor_bh30_264: Compressor_3_2
      port map ( R => CompressorOut_bh30_264_264,
                 X0 => CompressorIn_bh30_264_419);
   heap_bh30_w136_5 <= CompressorOut_bh30_264_264(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w137_6 <= CompressorOut_bh30_264_264(1); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_265_420 <= heap_bh30_w138_2 & heap_bh30_w138_1 & heap_bh30_w138_0;
      Compressor_bh30_265: Compressor_3_2
      port map ( R => CompressorOut_bh30_265_265,
                 X0 => CompressorIn_bh30_265_420);
   heap_bh30_w138_5 <= CompressorOut_bh30_265_265(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w139_6 <= CompressorOut_bh30_265_265(1); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_266_421 <= heap_bh30_w140_2 & heap_bh30_w140_1 & heap_bh30_w140_0;
      Compressor_bh30_266: Compressor_3_2
      port map ( R => CompressorOut_bh30_266_266,
                 X0 => CompressorIn_bh30_266_421);
   heap_bh30_w140_5 <= CompressorOut_bh30_266_266(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w141_6 <= CompressorOut_bh30_266_266(1); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_267_422 <= heap_bh30_w142_2 & heap_bh30_w142_1 & heap_bh30_w142_0;
      Compressor_bh30_267: Compressor_3_2
      port map ( R => CompressorOut_bh30_267_267,
                 X0 => CompressorIn_bh30_267_422);
   heap_bh30_w142_5 <= CompressorOut_bh30_267_267(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w143_6 <= CompressorOut_bh30_267_267(1); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_268_423 <= heap_bh30_w144_2 & heap_bh30_w144_1 & heap_bh30_w144_0;
      Compressor_bh30_268: Compressor_3_2
      port map ( R => CompressorOut_bh30_268_268,
                 X0 => CompressorIn_bh30_268_423);
   heap_bh30_w144_5 <= CompressorOut_bh30_268_268(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w145_6 <= CompressorOut_bh30_268_268(1); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_269_424 <= heap_bh30_w73_5 & heap_bh30_w73_4 & heap_bh30_w73_19 & heap_bh30_w73_18 & heap_bh30_w73_17 & heap_bh30_w73_16;
      Compressor_bh30_269: Compressor_6_3
      port map ( R => CompressorOut_bh30_269_269,
                 X0 => CompressorIn_bh30_269_424);
   heap_bh30_w73_20 <= CompressorOut_bh30_269_269(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w74_20 <= CompressorOut_bh30_269_269(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w75_21 <= CompressorOut_bh30_269_269(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_270_425 <= heap_bh30_w76_5 & heap_bh30_w76_4 & heap_bh30_w76_19 & heap_bh30_w76_18 & heap_bh30_w76_17 & heap_bh30_w76_16;
      Compressor_bh30_270: Compressor_6_3
      port map ( R => CompressorOut_bh30_270_270,
                 X0 => CompressorIn_bh30_270_425);
   heap_bh30_w76_20 <= CompressorOut_bh30_270_270(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w77_20 <= CompressorOut_bh30_270_270(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w78_21 <= CompressorOut_bh30_270_270(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_271_426 <= heap_bh30_w79_5 & heap_bh30_w79_4 & heap_bh30_w79_19 & heap_bh30_w79_18 & heap_bh30_w79_17 & heap_bh30_w79_16;
      Compressor_bh30_271: Compressor_6_3
      port map ( R => CompressorOut_bh30_271_271,
                 X0 => CompressorIn_bh30_271_426);
   heap_bh30_w79_20 <= CompressorOut_bh30_271_271(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w80_20 <= CompressorOut_bh30_271_271(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w81_21 <= CompressorOut_bh30_271_271(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_272_427 <= heap_bh30_w82_5 & heap_bh30_w82_4 & heap_bh30_w82_19 & heap_bh30_w82_18 & heap_bh30_w82_17 & heap_bh30_w82_16;
      Compressor_bh30_272: Compressor_6_3
      port map ( R => CompressorOut_bh30_272_272,
                 X0 => CompressorIn_bh30_272_427);
   heap_bh30_w82_20 <= CompressorOut_bh30_272_272(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w83_20 <= CompressorOut_bh30_272_272(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w84_21 <= CompressorOut_bh30_272_272(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_273_428 <= heap_bh30_w85_5 & heap_bh30_w85_4 & heap_bh30_w85_19 & heap_bh30_w85_18 & heap_bh30_w85_17 & heap_bh30_w85_16;
      Compressor_bh30_273: Compressor_6_3
      port map ( R => CompressorOut_bh30_273_273,
                 X0 => CompressorIn_bh30_273_428);
   heap_bh30_w85_20 <= CompressorOut_bh30_273_273(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w86_20 <= CompressorOut_bh30_273_273(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w87_21 <= CompressorOut_bh30_273_273(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_274_429 <= heap_bh30_w88_5 & heap_bh30_w88_4 & heap_bh30_w88_19 & heap_bh30_w88_18 & heap_bh30_w88_17 & heap_bh30_w88_16;
      Compressor_bh30_274: Compressor_6_3
      port map ( R => CompressorOut_bh30_274_274,
                 X0 => CompressorIn_bh30_274_429);
   heap_bh30_w88_20 <= CompressorOut_bh30_274_274(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w89_20 <= CompressorOut_bh30_274_274(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w90_20 <= CompressorOut_bh30_274_274(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_275_430 <= heap_bh30_w91_4 & heap_bh30_w91_3 & heap_bh30_w91_17 & heap_bh30_w91_16 & heap_bh30_w91_15 & heap_bh30_w91_14;
      Compressor_bh30_275: Compressor_6_3
      port map ( R => CompressorOut_bh30_275_275,
                 X0 => CompressorIn_bh30_275_430);
   heap_bh30_w91_18 <= CompressorOut_bh30_275_275(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w92_16 <= CompressorOut_bh30_275_275(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w93_15 <= CompressorOut_bh30_275_275(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_276_431 <= heap_bh30_w94_2 & heap_bh30_w94_1 & heap_bh30_w94_12 & heap_bh30_w94_11 & heap_bh30_w94_10 & heap_bh30_w94_9;
      Compressor_bh30_276: Compressor_6_3
      port map ( R => CompressorOut_bh30_276_276,
                 X0 => CompressorIn_bh30_276_431);
   heap_bh30_w94_13 <= CompressorOut_bh30_276_276(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w95_12 <= CompressorOut_bh30_276_276(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w96_11 <= CompressorOut_bh30_276_276(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_277_432 <= heap_bh30_w95_1 & heap_bh30_w95_0 & heap_bh30_w95_11 & heap_bh30_w95_10 & heap_bh30_w95_9 & heap_bh30_w95_8;
      Compressor_bh30_277: Compressor_6_3
      port map ( R => CompressorOut_bh30_277_277,
                 X0 => CompressorIn_bh30_277_432);
   heap_bh30_w95_13 <= CompressorOut_bh30_277_277(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w96_12 <= CompressorOut_bh30_277_277(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w97_11 <= CompressorOut_bh30_277_277(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_278_433 <= heap_bh30_w34_4 & heap_bh30_w34_14 & heap_bh30_w34_13 & heap_bh30_w34_12;
   CompressorIn_bh30_278_434(0) <= heap_bh30_w35_13;
      Compressor_bh30_278: Compressor_14_3
      port map ( R => CompressorOut_bh30_278_278,
                 X0 => CompressorIn_bh30_278_433,
                 X1 => CompressorIn_bh30_278_434);
   heap_bh30_w34_15 <= CompressorOut_bh30_278_278(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w35_14 <= CompressorOut_bh30_278_278(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w36_15 <= CompressorOut_bh30_278_278(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_279_435 <= heap_bh30_w37_4 & heap_bh30_w37_14 & heap_bh30_w37_13 & heap_bh30_w37_12;
   CompressorIn_bh30_279_436(0) <= heap_bh30_w38_13;
      Compressor_bh30_279: Compressor_14_3
      port map ( R => CompressorOut_bh30_279_279,
                 X0 => CompressorIn_bh30_279_435,
                 X1 => CompressorIn_bh30_279_436);
   heap_bh30_w37_15 <= CompressorOut_bh30_279_279(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w38_14 <= CompressorOut_bh30_279_279(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w39_15 <= CompressorOut_bh30_279_279(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_280_437 <= heap_bh30_w40_4 & heap_bh30_w40_14 & heap_bh30_w40_13 & heap_bh30_w40_12;
   CompressorIn_bh30_280_438(0) <= heap_bh30_w41_13;
      Compressor_bh30_280: Compressor_14_3
      port map ( R => CompressorOut_bh30_280_280,
                 X0 => CompressorIn_bh30_280_437,
                 X1 => CompressorIn_bh30_280_438);
   heap_bh30_w40_15 <= CompressorOut_bh30_280_280(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w41_14 <= CompressorOut_bh30_280_280(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w42_15 <= CompressorOut_bh30_280_280(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_281_439 <= heap_bh30_w43_4 & heap_bh30_w43_14 & heap_bh30_w43_13 & heap_bh30_w43_12;
   CompressorIn_bh30_281_440(0) <= heap_bh30_w44_13;
      Compressor_bh30_281: Compressor_14_3
      port map ( R => CompressorOut_bh30_281_281,
                 X0 => CompressorIn_bh30_281_439,
                 X1 => CompressorIn_bh30_281_440);
   heap_bh30_w43_15 <= CompressorOut_bh30_281_281(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w44_14 <= CompressorOut_bh30_281_281(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w45_15 <= CompressorOut_bh30_281_281(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_282_441 <= heap_bh30_w48_4 & heap_bh30_w48_15 & heap_bh30_w48_14 & heap_bh30_w48_13;
   CompressorIn_bh30_282_442(0) <= heap_bh30_w49_15;
      Compressor_bh30_282: Compressor_14_3
      port map ( R => CompressorOut_bh30_282_282,
                 X0 => CompressorIn_bh30_282_441,
                 X1 => CompressorIn_bh30_282_442);
   heap_bh30_w48_16 <= CompressorOut_bh30_282_282(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w49_16 <= CompressorOut_bh30_282_282(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w50_16 <= CompressorOut_bh30_282_282(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_283_443 <= heap_bh30_w50_3 & heap_bh30_w50_15 & heap_bh30_w50_14 & heap_bh30_w50_13;
   CompressorIn_bh30_283_444(0) <= heap_bh30_w51_5;
      Compressor_bh30_283: Compressor_14_3
      port map ( R => CompressorOut_bh30_283_283,
                 X0 => CompressorIn_bh30_283_443,
                 X1 => CompressorIn_bh30_283_444);
   heap_bh30_w50_17 <= CompressorOut_bh30_283_283(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w51_17 <= CompressorOut_bh30_283_283(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w52_17 <= CompressorOut_bh30_283_283(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_284_445 <= heap_bh30_w51_4 & heap_bh30_w51_16 & heap_bh30_w51_15 & heap_bh30_w51_14;
   CompressorIn_bh30_284_446(0) <= heap_bh30_w52_4;
      Compressor_bh30_284: Compressor_14_3
      port map ( R => CompressorOut_bh30_284_284,
                 X0 => CompressorIn_bh30_284_445,
                 X1 => CompressorIn_bh30_284_446);
   heap_bh30_w51_18 <= CompressorOut_bh30_284_284(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w52_18 <= CompressorOut_bh30_284_284(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w53_16 <= CompressorOut_bh30_284_284(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_285_447 <= heap_bh30_w53_3 & heap_bh30_w53_15 & heap_bh30_w53_14 & heap_bh30_w53_13;
   CompressorIn_bh30_285_448(0) <= heap_bh30_w54_5;
      Compressor_bh30_285: Compressor_14_3
      port map ( R => CompressorOut_bh30_285_285,
                 X0 => CompressorIn_bh30_285_447,
                 X1 => CompressorIn_bh30_285_448);
   heap_bh30_w53_17 <= CompressorOut_bh30_285_285(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w54_17 <= CompressorOut_bh30_285_285(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w55_17 <= CompressorOut_bh30_285_285(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_286_449 <= heap_bh30_w54_4 & heap_bh30_w54_16 & heap_bh30_w54_15 & heap_bh30_w54_14;
   CompressorIn_bh30_286_450(0) <= heap_bh30_w55_4;
      Compressor_bh30_286: Compressor_14_3
      port map ( R => CompressorOut_bh30_286_286,
                 X0 => CompressorIn_bh30_286_449,
                 X1 => CompressorIn_bh30_286_450);
   heap_bh30_w54_18 <= CompressorOut_bh30_286_286(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w55_18 <= CompressorOut_bh30_286_286(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w56_16 <= CompressorOut_bh30_286_286(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_287_451 <= heap_bh30_w56_3 & heap_bh30_w56_15 & heap_bh30_w56_14 & heap_bh30_w56_13;
   CompressorIn_bh30_287_452(0) <= heap_bh30_w57_5;
      Compressor_bh30_287: Compressor_14_3
      port map ( R => CompressorOut_bh30_287_287,
                 X0 => CompressorIn_bh30_287_451,
                 X1 => CompressorIn_bh30_287_452);
   heap_bh30_w56_17 <= CompressorOut_bh30_287_287(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w57_17 <= CompressorOut_bh30_287_287(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w58_17 <= CompressorOut_bh30_287_287(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_288_453 <= heap_bh30_w57_4 & heap_bh30_w57_16 & heap_bh30_w57_15 & heap_bh30_w57_14;
   CompressorIn_bh30_288_454(0) <= heap_bh30_w58_4;
      Compressor_bh30_288: Compressor_14_3
      port map ( R => CompressorOut_bh30_288_288,
                 X0 => CompressorIn_bh30_288_453,
                 X1 => CompressorIn_bh30_288_454);
   heap_bh30_w57_18 <= CompressorOut_bh30_288_288(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w58_18 <= CompressorOut_bh30_288_288(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w59_16 <= CompressorOut_bh30_288_288(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_289_455 <= heap_bh30_w59_3 & heap_bh30_w59_15 & heap_bh30_w59_14 & heap_bh30_w59_13;
   CompressorIn_bh30_289_456(0) <= heap_bh30_w60_5;
      Compressor_bh30_289: Compressor_14_3
      port map ( R => CompressorOut_bh30_289_289,
                 X0 => CompressorIn_bh30_289_455,
                 X1 => CompressorIn_bh30_289_456);
   heap_bh30_w59_17 <= CompressorOut_bh30_289_289(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w60_17 <= CompressorOut_bh30_289_289(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w61_17 <= CompressorOut_bh30_289_289(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_290_457 <= heap_bh30_w60_4 & heap_bh30_w60_16 & heap_bh30_w60_15 & heap_bh30_w60_14;
   CompressorIn_bh30_290_458(0) <= heap_bh30_w61_4;
      Compressor_bh30_290: Compressor_14_3
      port map ( R => CompressorOut_bh30_290_290,
                 X0 => CompressorIn_bh30_290_457,
                 X1 => CompressorIn_bh30_290_458);
   heap_bh30_w60_18 <= CompressorOut_bh30_290_290(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w61_18 <= CompressorOut_bh30_290_290(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w62_16 <= CompressorOut_bh30_290_290(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_291_459 <= heap_bh30_w62_3 & heap_bh30_w62_15 & heap_bh30_w62_14 & heap_bh30_w62_13;
   CompressorIn_bh30_291_460(0) <= heap_bh30_w63_5;
      Compressor_bh30_291: Compressor_14_3
      port map ( R => CompressorOut_bh30_291_291,
                 X0 => CompressorIn_bh30_291_459,
                 X1 => CompressorIn_bh30_291_460);
   heap_bh30_w62_17 <= CompressorOut_bh30_291_291(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w63_17 <= CompressorOut_bh30_291_291(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w64_17 <= CompressorOut_bh30_291_291(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_292_461 <= heap_bh30_w63_4 & heap_bh30_w63_16 & heap_bh30_w63_15 & heap_bh30_w63_14;
   CompressorIn_bh30_292_462(0) <= heap_bh30_w64_4;
      Compressor_bh30_292: Compressor_14_3
      port map ( R => CompressorOut_bh30_292_292,
                 X0 => CompressorIn_bh30_292_461,
                 X1 => CompressorIn_bh30_292_462);
   heap_bh30_w63_18 <= CompressorOut_bh30_292_292(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w64_18 <= CompressorOut_bh30_292_292(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w65_16 <= CompressorOut_bh30_292_292(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_293_463 <= heap_bh30_w65_3 & heap_bh30_w65_15 & heap_bh30_w65_14 & heap_bh30_w65_13;
   CompressorIn_bh30_293_464(0) <= heap_bh30_w66_5;
      Compressor_bh30_293: Compressor_14_3
      port map ( R => CompressorOut_bh30_293_293,
                 X0 => CompressorIn_bh30_293_463,
                 X1 => CompressorIn_bh30_293_464);
   heap_bh30_w65_17 <= CompressorOut_bh30_293_293(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w66_17 <= CompressorOut_bh30_293_293(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w67_18 <= CompressorOut_bh30_293_293(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_294_465 <= heap_bh30_w66_4 & heap_bh30_w66_16 & heap_bh30_w66_15 & heap_bh30_w66_14;
   CompressorIn_bh30_294_466(0) <= heap_bh30_w67_5;
      Compressor_bh30_294: Compressor_14_3
      port map ( R => CompressorOut_bh30_294_294,
                 X0 => CompressorIn_bh30_294_465,
                 X1 => CompressorIn_bh30_294_466);
   heap_bh30_w66_18 <= CompressorOut_bh30_294_294(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w67_19 <= CompressorOut_bh30_294_294(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w68_17 <= CompressorOut_bh30_294_294(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_295_467 <= heap_bh30_w67_4 & heap_bh30_w67_17 & heap_bh30_w67_16 & heap_bh30_w67_15;
   CompressorIn_bh30_295_468(0) <= heap_bh30_w68_4;
      Compressor_bh30_295: Compressor_14_3
      port map ( R => CompressorOut_bh30_295_295,
                 X0 => CompressorIn_bh30_295_467,
                 X1 => CompressorIn_bh30_295_468);
   heap_bh30_w67_20 <= CompressorOut_bh30_295_295(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w68_18 <= CompressorOut_bh30_295_295(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w69_19 <= CompressorOut_bh30_295_295(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_296_469 <= heap_bh30_w68_3 & heap_bh30_w68_16 & heap_bh30_w68_15 & heap_bh30_w68_14;
   CompressorIn_bh30_296_470(0) <= heap_bh30_w69_18;
      Compressor_bh30_296: Compressor_14_3
      port map ( R => CompressorOut_bh30_296_296,
                 X0 => CompressorIn_bh30_296_469,
                 X1 => CompressorIn_bh30_296_470);
   heap_bh30_w68_19 <= CompressorOut_bh30_296_296(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w69_20 <= CompressorOut_bh30_296_296(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w70_19 <= CompressorOut_bh30_296_296(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_297_471 <= heap_bh30_w70_18 & heap_bh30_w70_17 & heap_bh30_w70_16 & heap_bh30_w70_15;
   CompressorIn_bh30_297_472(0) <= heap_bh30_w71_19;
      Compressor_bh30_297: Compressor_14_3
      port map ( R => CompressorOut_bh30_297_297,
                 X0 => CompressorIn_bh30_297_471,
                 X1 => CompressorIn_bh30_297_472);
   heap_bh30_w70_20 <= CompressorOut_bh30_297_297(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w71_20 <= CompressorOut_bh30_297_297(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w72_21 <= CompressorOut_bh30_297_297(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_298_473 <= heap_bh30_w71_18 & heap_bh30_w71_17 & heap_bh30_w71_16 & heap_bh30_w71_15;
   CompressorIn_bh30_298_474(0) <= heap_bh30_w72_20;
      Compressor_bh30_298: Compressor_14_3
      port map ( R => CompressorOut_bh30_298_298,
                 X0 => CompressorIn_bh30_298_473,
                 X1 => CompressorIn_bh30_298_474);
   heap_bh30_w71_21 <= CompressorOut_bh30_298_298(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w72_22 <= CompressorOut_bh30_298_298(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w73_21 <= CompressorOut_bh30_298_298(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_299_475 <= heap_bh30_w74_19 & heap_bh30_w74_18 & heap_bh30_w74_17 & heap_bh30_w74_16;
   CompressorIn_bh30_299_476(0) <= heap_bh30_w75_20;
      Compressor_bh30_299: Compressor_14_3
      port map ( R => CompressorOut_bh30_299_299,
                 X0 => CompressorIn_bh30_299_475,
                 X1 => CompressorIn_bh30_299_476);
   heap_bh30_w74_21 <= CompressorOut_bh30_299_299(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w75_22 <= CompressorOut_bh30_299_299(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w76_21 <= CompressorOut_bh30_299_299(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_300_477 <= heap_bh30_w77_19 & heap_bh30_w77_18 & heap_bh30_w77_17 & heap_bh30_w77_16;
   CompressorIn_bh30_300_478(0) <= heap_bh30_w78_20;
      Compressor_bh30_300: Compressor_14_3
      port map ( R => CompressorOut_bh30_300_300,
                 X0 => CompressorIn_bh30_300_477,
                 X1 => CompressorIn_bh30_300_478);
   heap_bh30_w77_21 <= CompressorOut_bh30_300_300(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w78_22 <= CompressorOut_bh30_300_300(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w79_21 <= CompressorOut_bh30_300_300(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_301_479 <= heap_bh30_w80_19 & heap_bh30_w80_18 & heap_bh30_w80_17 & heap_bh30_w80_16;
   CompressorIn_bh30_301_480(0) <= heap_bh30_w81_20;
      Compressor_bh30_301: Compressor_14_3
      port map ( R => CompressorOut_bh30_301_301,
                 X0 => CompressorIn_bh30_301_479,
                 X1 => CompressorIn_bh30_301_480);
   heap_bh30_w80_21 <= CompressorOut_bh30_301_301(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w81_22 <= CompressorOut_bh30_301_301(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w82_21 <= CompressorOut_bh30_301_301(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_302_481 <= heap_bh30_w83_19 & heap_bh30_w83_18 & heap_bh30_w83_17 & heap_bh30_w83_16;
   CompressorIn_bh30_302_482(0) <= heap_bh30_w84_20;
      Compressor_bh30_302: Compressor_14_3
      port map ( R => CompressorOut_bh30_302_302,
                 X0 => CompressorIn_bh30_302_481,
                 X1 => CompressorIn_bh30_302_482);
   heap_bh30_w83_21 <= CompressorOut_bh30_302_302(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w84_22 <= CompressorOut_bh30_302_302(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w85_21 <= CompressorOut_bh30_302_302(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_303_483 <= heap_bh30_w86_19 & heap_bh30_w86_18 & heap_bh30_w86_17 & heap_bh30_w86_16;
   CompressorIn_bh30_303_484(0) <= heap_bh30_w87_20;
      Compressor_bh30_303: Compressor_14_3
      port map ( R => CompressorOut_bh30_303_303,
                 X0 => CompressorIn_bh30_303_483,
                 X1 => CompressorIn_bh30_303_484);
   heap_bh30_w86_21 <= CompressorOut_bh30_303_303(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w87_22 <= CompressorOut_bh30_303_303(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w88_21 <= CompressorOut_bh30_303_303(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_304_485 <= heap_bh30_w89_19 & heap_bh30_w89_18 & heap_bh30_w89_17 & heap_bh30_w89_16;
   CompressorIn_bh30_304_486(0) <= heap_bh30_w90_19;
      Compressor_bh30_304: Compressor_14_3
      port map ( R => CompressorOut_bh30_304_304,
                 X0 => CompressorIn_bh30_304_485,
                 X1 => CompressorIn_bh30_304_486);
   heap_bh30_w89_21 <= CompressorOut_bh30_304_304(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w90_21 <= CompressorOut_bh30_304_304(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w91_19 <= CompressorOut_bh30_304_304(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_305_487 <= heap_bh30_w92_15 & heap_bh30_w92_14 & heap_bh30_w92_13 & heap_bh30_w92_12;
   CompressorIn_bh30_305_488(0) <= heap_bh30_w93_14;
      Compressor_bh30_305: Compressor_14_3
      port map ( R => CompressorOut_bh30_305_305,
                 X0 => CompressorIn_bh30_305_487,
                 X1 => CompressorIn_bh30_305_488);
   heap_bh30_w92_17 <= CompressorOut_bh30_305_305(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w93_16 <= CompressorOut_bh30_305_305(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w94_14 <= CompressorOut_bh30_305_305(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_306_489 <= heap_bh30_w96_1 & heap_bh30_w96_0 & heap_bh30_w96_10 & heap_bh30_w96_9;
   CompressorIn_bh30_306_490(0) <= heap_bh30_w97_1;
      Compressor_bh30_306: Compressor_14_3
      port map ( R => CompressorOut_bh30_306_306,
                 X0 => CompressorIn_bh30_306_489,
                 X1 => CompressorIn_bh30_306_490);
   heap_bh30_w96_13 <= CompressorOut_bh30_306_306(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w97_12 <= CompressorOut_bh30_306_306(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w98_11 <= CompressorOut_bh30_306_306(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_307_491 <= heap_bh30_w97_0 & heap_bh30_w97_10 & heap_bh30_w97_9 & heap_bh30_w97_8;
   CompressorIn_bh30_307_492(0) <= heap_bh30_w98_1;
      Compressor_bh30_307: Compressor_14_3
      port map ( R => CompressorOut_bh30_307_307,
                 X0 => CompressorIn_bh30_307_491,
                 X1 => CompressorIn_bh30_307_492);
   heap_bh30_w97_13 <= CompressorOut_bh30_307_307(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w98_12 <= CompressorOut_bh30_307_307(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w99_11 <= CompressorOut_bh30_307_307(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_308_493 <= heap_bh30_w98_0 & heap_bh30_w98_10 & heap_bh30_w98_9 & heap_bh30_w98_8;
   CompressorIn_bh30_308_494(0) <= heap_bh30_w99_1;
      Compressor_bh30_308: Compressor_14_3
      port map ( R => CompressorOut_bh30_308_308,
                 X0 => CompressorIn_bh30_308_493,
                 X1 => CompressorIn_bh30_308_494);
   heap_bh30_w98_13 <= CompressorOut_bh30_308_308(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w99_12 <= CompressorOut_bh30_308_308(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w100_11 <= CompressorOut_bh30_308_308(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_309_495 <= heap_bh30_w99_0 & heap_bh30_w99_10 & heap_bh30_w99_9 & heap_bh30_w99_8;
   CompressorIn_bh30_309_496(0) <= heap_bh30_w100_1;
      Compressor_bh30_309: Compressor_14_3
      port map ( R => CompressorOut_bh30_309_309,
                 X0 => CompressorIn_bh30_309_495,
                 X1 => CompressorIn_bh30_309_496);
   heap_bh30_w99_13 <= CompressorOut_bh30_309_309(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w100_12 <= CompressorOut_bh30_309_309(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w101_11 <= CompressorOut_bh30_309_309(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_310_497 <= heap_bh30_w100_0 & heap_bh30_w100_10 & heap_bh30_w100_9 & heap_bh30_w100_8;
   CompressorIn_bh30_310_498(0) <= heap_bh30_w101_1;
      Compressor_bh30_310: Compressor_14_3
      port map ( R => CompressorOut_bh30_310_310,
                 X0 => CompressorIn_bh30_310_497,
                 X1 => CompressorIn_bh30_310_498);
   heap_bh30_w100_13 <= CompressorOut_bh30_310_310(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w101_12 <= CompressorOut_bh30_310_310(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w102_11 <= CompressorOut_bh30_310_310(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_311_499 <= heap_bh30_w101_0 & heap_bh30_w101_10 & heap_bh30_w101_9 & heap_bh30_w101_8;
   CompressorIn_bh30_311_500(0) <= heap_bh30_w102_1;
      Compressor_bh30_311: Compressor_14_3
      port map ( R => CompressorOut_bh30_311_311,
                 X0 => CompressorIn_bh30_311_499,
                 X1 => CompressorIn_bh30_311_500);
   heap_bh30_w101_13 <= CompressorOut_bh30_311_311(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w102_12 <= CompressorOut_bh30_311_311(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w103_11 <= CompressorOut_bh30_311_311(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_312_501 <= heap_bh30_w102_0 & heap_bh30_w102_10 & heap_bh30_w102_9 & heap_bh30_w102_8;
   CompressorIn_bh30_312_502(0) <= heap_bh30_w103_1;
      Compressor_bh30_312: Compressor_14_3
      port map ( R => CompressorOut_bh30_312_312,
                 X0 => CompressorIn_bh30_312_501,
                 X1 => CompressorIn_bh30_312_502);
   heap_bh30_w102_13 <= CompressorOut_bh30_312_312(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w103_12 <= CompressorOut_bh30_312_312(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w104_11 <= CompressorOut_bh30_312_312(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_313_503 <= heap_bh30_w103_0 & heap_bh30_w103_10 & heap_bh30_w103_9 & heap_bh30_w103_8;
   CompressorIn_bh30_313_504(0) <= heap_bh30_w104_1;
      Compressor_bh30_313: Compressor_14_3
      port map ( R => CompressorOut_bh30_313_313,
                 X0 => CompressorIn_bh30_313_503,
                 X1 => CompressorIn_bh30_313_504);
   heap_bh30_w103_13 <= CompressorOut_bh30_313_313(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w104_12 <= CompressorOut_bh30_313_313(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w105_11 <= CompressorOut_bh30_313_313(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_314_505 <= heap_bh30_w104_0 & heap_bh30_w104_10 & heap_bh30_w104_9 & heap_bh30_w104_8;
   CompressorIn_bh30_314_506(0) <= heap_bh30_w105_1;
      Compressor_bh30_314: Compressor_14_3
      port map ( R => CompressorOut_bh30_314_314,
                 X0 => CompressorIn_bh30_314_505,
                 X1 => CompressorIn_bh30_314_506);
   heap_bh30_w104_13 <= CompressorOut_bh30_314_314(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w105_12 <= CompressorOut_bh30_314_314(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w106_11 <= CompressorOut_bh30_314_314(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_315_507 <= heap_bh30_w105_0 & heap_bh30_w105_10 & heap_bh30_w105_9 & heap_bh30_w105_8;
   CompressorIn_bh30_315_508(0) <= heap_bh30_w106_1;
      Compressor_bh30_315: Compressor_14_3
      port map ( R => CompressorOut_bh30_315_315,
                 X0 => CompressorIn_bh30_315_507,
                 X1 => CompressorIn_bh30_315_508);
   heap_bh30_w105_13 <= CompressorOut_bh30_315_315(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w106_12 <= CompressorOut_bh30_315_315(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w107_11 <= CompressorOut_bh30_315_315(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_316_509 <= heap_bh30_w106_0 & heap_bh30_w106_10 & heap_bh30_w106_9 & heap_bh30_w106_8;
   CompressorIn_bh30_316_510(0) <= heap_bh30_w107_1;
      Compressor_bh30_316: Compressor_14_3
      port map ( R => CompressorOut_bh30_316_316,
                 X0 => CompressorIn_bh30_316_509,
                 X1 => CompressorIn_bh30_316_510);
   heap_bh30_w106_13 <= CompressorOut_bh30_316_316(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w107_12 <= CompressorOut_bh30_316_316(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w108_10 <= CompressorOut_bh30_316_316(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_317_511 <= heap_bh30_w107_0 & heap_bh30_w107_10 & heap_bh30_w107_9 & heap_bh30_w107_8;
   CompressorIn_bh30_317_512(0) <= heap_bh30_w108_0;
      Compressor_bh30_317: Compressor_14_3
      port map ( R => CompressorOut_bh30_317_317,
                 X0 => CompressorIn_bh30_317_511,
                 X1 => CompressorIn_bh30_317_512);
   heap_bh30_w107_13 <= CompressorOut_bh30_317_317(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w108_11 <= CompressorOut_bh30_317_317(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w109_10 <= CompressorOut_bh30_317_317(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_318_513 <= heap_bh30_w109_0 & heap_bh30_w109_9 & heap_bh30_w109_8 & heap_bh30_w109_7;
   CompressorIn_bh30_318_514(0) <= heap_bh30_w110_0;
      Compressor_bh30_318: Compressor_14_3
      port map ( R => CompressorOut_bh30_318_318,
                 X0 => CompressorIn_bh30_318_513,
                 X1 => CompressorIn_bh30_318_514);
   heap_bh30_w109_11 <= CompressorOut_bh30_318_318(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w110_10 <= CompressorOut_bh30_318_318(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w111_10 <= CompressorOut_bh30_318_318(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_319_515 <= heap_bh30_w111_0 & heap_bh30_w111_9 & heap_bh30_w111_8 & heap_bh30_w111_7;
   CompressorIn_bh30_319_516(0) <= heap_bh30_w112_8;
      Compressor_bh30_319: Compressor_14_3
      port map ( R => CompressorOut_bh30_319_319,
                 X0 => CompressorIn_bh30_319_515,
                 X1 => CompressorIn_bh30_319_516);
   heap_bh30_w111_11 <= CompressorOut_bh30_319_319(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w112_9 <= CompressorOut_bh30_319_319(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w113_9 <= CompressorOut_bh30_319_319(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_320_517 <= heap_bh30_w129_0 & heap_bh30_w129_7 & heap_bh30_w129_6 & heap_bh30_w129_5;
   CompressorIn_bh30_320_518(0) <= heap_bh30_w130_7;
      Compressor_bh30_320: Compressor_14_3
      port map ( R => CompressorOut_bh30_320_320,
                 X0 => CompressorIn_bh30_320_517,
                 X1 => CompressorIn_bh30_320_518);
   heap_bh30_w129_8 <= CompressorOut_bh30_320_320(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w130_8 <= CompressorOut_bh30_320_320(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w131_8 <= CompressorOut_bh30_320_320(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_321_519 <= heap_bh30_w72_19 & heap_bh30_w72_18 & heap_bh30_w72_17 & heap_bh30_w72_16;
      Compressor_bh30_321: Compressor_4_3
      port map ( R => CompressorOut_bh30_321_321,
                 X0 => CompressorIn_bh30_321_519);
   heap_bh30_w72_23 <= CompressorOut_bh30_321_321(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w73_22 <= CompressorOut_bh30_321_321(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w74_22 <= CompressorOut_bh30_321_321(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_322_520 <= heap_bh30_w75_19 & heap_bh30_w75_18 & heap_bh30_w75_17 & heap_bh30_w75_16;
      Compressor_bh30_322: Compressor_4_3
      port map ( R => CompressorOut_bh30_322_322,
                 X0 => CompressorIn_bh30_322_520);
   heap_bh30_w75_23 <= CompressorOut_bh30_322_322(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w76_22 <= CompressorOut_bh30_322_322(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w77_22 <= CompressorOut_bh30_322_322(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_323_521 <= heap_bh30_w78_19 & heap_bh30_w78_18 & heap_bh30_w78_17 & heap_bh30_w78_16;
      Compressor_bh30_323: Compressor_4_3
      port map ( R => CompressorOut_bh30_323_323,
                 X0 => CompressorIn_bh30_323_521);
   heap_bh30_w78_23 <= CompressorOut_bh30_323_323(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w79_22 <= CompressorOut_bh30_323_323(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w80_22 <= CompressorOut_bh30_323_323(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_324_522 <= heap_bh30_w81_19 & heap_bh30_w81_18 & heap_bh30_w81_17 & heap_bh30_w81_16;
      Compressor_bh30_324: Compressor_4_3
      port map ( R => CompressorOut_bh30_324_324,
                 X0 => CompressorIn_bh30_324_522);
   heap_bh30_w81_23 <= CompressorOut_bh30_324_324(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w82_22 <= CompressorOut_bh30_324_324(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w83_22 <= CompressorOut_bh30_324_324(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_325_523 <= heap_bh30_w84_19 & heap_bh30_w84_18 & heap_bh30_w84_17 & heap_bh30_w84_16;
      Compressor_bh30_325: Compressor_4_3
      port map ( R => CompressorOut_bh30_325_325,
                 X0 => CompressorIn_bh30_325_523);
   heap_bh30_w84_23 <= CompressorOut_bh30_325_325(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w85_22 <= CompressorOut_bh30_325_325(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w86_22 <= CompressorOut_bh30_325_325(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_326_524 <= heap_bh30_w87_19 & heap_bh30_w87_18 & heap_bh30_w87_17 & heap_bh30_w87_16;
      Compressor_bh30_326: Compressor_4_3
      port map ( R => CompressorOut_bh30_326_326,
                 X0 => CompressorIn_bh30_326_524);
   heap_bh30_w87_23 <= CompressorOut_bh30_326_326(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w88_22 <= CompressorOut_bh30_326_326(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w89_22 <= CompressorOut_bh30_326_326(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_327_525 <= heap_bh30_w90_18 & heap_bh30_w90_17 & heap_bh30_w90_16 & heap_bh30_w90_15;
      Compressor_bh30_327: Compressor_4_3
      port map ( R => CompressorOut_bh30_327_327,
                 X0 => CompressorIn_bh30_327_525);
   heap_bh30_w90_22 <= CompressorOut_bh30_327_327(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w91_20 <= CompressorOut_bh30_327_327(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w92_18 <= CompressorOut_bh30_327_327(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_328_526 <= heap_bh30_w93_13 & heap_bh30_w93_12 & heap_bh30_w93_11 & heap_bh30_w93_10;
      Compressor_bh30_328: Compressor_4_3
      port map ( R => CompressorOut_bh30_328_328,
                 X0 => CompressorIn_bh30_328_526);
   heap_bh30_w93_17 <= CompressorOut_bh30_328_328(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w94_15 <= CompressorOut_bh30_328_328(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w95_14 <= CompressorOut_bh30_328_328(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_329_527 <= heap_bh30_w8_6 & heap_bh30_w8_3 & heap_bh30_w8_7;
   CompressorIn_bh30_329_528 <= heap_bh30_w9_7 & heap_bh30_w9_4;
      Compressor_bh30_329: Compressor_23_3
      port map ( R => CompressorOut_bh30_329_329,
                 X0 => CompressorIn_bh30_329_527,
                 X1 => CompressorIn_bh30_329_528);
   heap_bh30_w8_8 <= CompressorOut_bh30_329_329(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w9_8 <= CompressorOut_bh30_329_329(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w10_9 <= CompressorOut_bh30_329_329(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_330_529 <= heap_bh30_w19_5 & heap_bh30_w19_4 & heap_bh30_w19_10;
   CompressorIn_bh30_330_530 <= heap_bh30_w20_10 & heap_bh30_w20_9;
      Compressor_bh30_330: Compressor_23_3
      port map ( R => CompressorOut_bh30_330_330,
                 X0 => CompressorIn_bh30_330_529,
                 X1 => CompressorIn_bh30_330_530);
   heap_bh30_w19_11 <= CompressorOut_bh30_330_330(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w20_11 <= CompressorOut_bh30_330_330(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w21_12 <= CompressorOut_bh30_330_330(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_331_531 <= heap_bh30_w22_5 & heap_bh30_w22_4 & heap_bh30_w22_10;
   CompressorIn_bh30_331_532 <= heap_bh30_w23_11 & heap_bh30_w23_10;
      Compressor_bh30_331: Compressor_23_3
      port map ( R => CompressorOut_bh30_331_331,
                 X0 => CompressorIn_bh30_331_531,
                 X1 => CompressorIn_bh30_331_532);
   heap_bh30_w22_11 <= CompressorOut_bh30_331_331(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w23_12 <= CompressorOut_bh30_331_331(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w24_13 <= CompressorOut_bh30_331_331(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_332_533 <= heap_bh30_w25_13 & heap_bh30_w25_12 & heap_bh30_w25_11;
   CompressorIn_bh30_332_534 <= heap_bh30_w26_12 & heap_bh30_w26_11;
      Compressor_bh30_332: Compressor_23_3
      port map ( R => CompressorOut_bh30_332_332,
                 X0 => CompressorIn_bh30_332_533,
                 X1 => CompressorIn_bh30_332_534);
   heap_bh30_w25_14 <= CompressorOut_bh30_332_332(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w26_13 <= CompressorOut_bh30_332_332(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w27_13 <= CompressorOut_bh30_332_332(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_333_535 <= heap_bh30_w28_13 & heap_bh30_w28_12 & heap_bh30_w28_11;
   CompressorIn_bh30_333_536 <= heap_bh30_w29_12 & heap_bh30_w29_11;
      Compressor_bh30_333: Compressor_23_3
      port map ( R => CompressorOut_bh30_333_333,
                 X0 => CompressorIn_bh30_333_535,
                 X1 => CompressorIn_bh30_333_536);
   heap_bh30_w28_14 <= CompressorOut_bh30_333_333(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w29_13 <= CompressorOut_bh30_333_333(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w30_13 <= CompressorOut_bh30_333_333(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_334_537 <= heap_bh30_w31_13 & heap_bh30_w31_12 & heap_bh30_w31_11;
   CompressorIn_bh30_334_538 <= heap_bh30_w32_12 & heap_bh30_w32_11;
      Compressor_bh30_334: Compressor_23_3
      port map ( R => CompressorOut_bh30_334_334,
                 X0 => CompressorIn_bh30_334_537,
                 X1 => CompressorIn_bh30_334_538);
   heap_bh30_w31_14 <= CompressorOut_bh30_334_334(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w32_13 <= CompressorOut_bh30_334_334(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w33_14 <= CompressorOut_bh30_334_334(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_335_539 <= heap_bh30_w45_14 & heap_bh30_w45_13 & heap_bh30_w45_12;
   CompressorIn_bh30_335_540 <= heap_bh30_w46_14 & heap_bh30_w46_13;
      Compressor_bh30_335: Compressor_23_3
      port map ( R => CompressorOut_bh30_335_335,
                 X0 => CompressorIn_bh30_335_539,
                 X1 => CompressorIn_bh30_335_540);
   heap_bh30_w45_16 <= CompressorOut_bh30_335_335(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w46_15 <= CompressorOut_bh30_335_335(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w47_15 <= CompressorOut_bh30_335_335(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_336_541 <= heap_bh30_w113_8 & heap_bh30_w113_7 & heap_bh30_w113_6;
   CompressorIn_bh30_336_542 <= heap_bh30_w114_8 & heap_bh30_w114_7;
      Compressor_bh30_336: Compressor_23_3
      port map ( R => CompressorOut_bh30_336_336,
                 X0 => CompressorIn_bh30_336_541,
                 X1 => CompressorIn_bh30_336_542);
   heap_bh30_w113_10 <= CompressorOut_bh30_336_336(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w114_9 <= CompressorOut_bh30_336_336(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w115_9 <= CompressorOut_bh30_336_336(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_337_543 <= heap_bh30_w115_8 & heap_bh30_w115_7 & heap_bh30_w115_6;
   CompressorIn_bh30_337_544 <= heap_bh30_w116_8 & heap_bh30_w116_7;
      Compressor_bh30_337: Compressor_23_3
      port map ( R => CompressorOut_bh30_337_337,
                 X0 => CompressorIn_bh30_337_543,
                 X1 => CompressorIn_bh30_337_544);
   heap_bh30_w115_10 <= CompressorOut_bh30_337_337(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w116_9 <= CompressorOut_bh30_337_337(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w117_9 <= CompressorOut_bh30_337_337(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_338_545 <= heap_bh30_w117_8 & heap_bh30_w117_7 & heap_bh30_w117_6;
   CompressorIn_bh30_338_546 <= heap_bh30_w118_8 & heap_bh30_w118_7;
      Compressor_bh30_338: Compressor_23_3
      port map ( R => CompressorOut_bh30_338_338,
                 X0 => CompressorIn_bh30_338_545,
                 X1 => CompressorIn_bh30_338_546);
   heap_bh30_w117_10 <= CompressorOut_bh30_338_338(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w118_9 <= CompressorOut_bh30_338_338(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w119_9 <= CompressorOut_bh30_338_338(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_339_547 <= heap_bh30_w119_8 & heap_bh30_w119_7 & heap_bh30_w119_6;
   CompressorIn_bh30_339_548 <= heap_bh30_w120_8 & heap_bh30_w120_7;
      Compressor_bh30_339: Compressor_23_3
      port map ( R => CompressorOut_bh30_339_339,
                 X0 => CompressorIn_bh30_339_547,
                 X1 => CompressorIn_bh30_339_548);
   heap_bh30_w119_10 <= CompressorOut_bh30_339_339(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w120_9 <= CompressorOut_bh30_339_339(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w121_9 <= CompressorOut_bh30_339_339(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_340_549 <= heap_bh30_w121_8 & heap_bh30_w121_7 & heap_bh30_w121_6;
   CompressorIn_bh30_340_550 <= heap_bh30_w122_8 & heap_bh30_w122_7;
      Compressor_bh30_340: Compressor_23_3
      port map ( R => CompressorOut_bh30_340_340,
                 X0 => CompressorIn_bh30_340_549,
                 X1 => CompressorIn_bh30_340_550);
   heap_bh30_w121_10 <= CompressorOut_bh30_340_340(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w122_9 <= CompressorOut_bh30_340_340(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w123_9 <= CompressorOut_bh30_340_340(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_341_551 <= heap_bh30_w123_8 & heap_bh30_w123_7 & heap_bh30_w123_6;
   CompressorIn_bh30_341_552 <= heap_bh30_w124_8 & heap_bh30_w124_7;
      Compressor_bh30_341: Compressor_23_3
      port map ( R => CompressorOut_bh30_341_341,
                 X0 => CompressorIn_bh30_341_551,
                 X1 => CompressorIn_bh30_341_552);
   heap_bh30_w123_10 <= CompressorOut_bh30_341_341(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w124_9 <= CompressorOut_bh30_341_341(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w125_9 <= CompressorOut_bh30_341_341(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_342_553 <= heap_bh30_w125_8 & heap_bh30_w125_7 & heap_bh30_w125_6;
   CompressorIn_bh30_342_554 <= heap_bh30_w126_8 & heap_bh30_w126_7;
      Compressor_bh30_342: Compressor_23_3
      port map ( R => CompressorOut_bh30_342_342,
                 X0 => CompressorIn_bh30_342_553,
                 X1 => CompressorIn_bh30_342_554);
   heap_bh30_w125_10 <= CompressorOut_bh30_342_342(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w126_9 <= CompressorOut_bh30_342_342(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w127_9 <= CompressorOut_bh30_342_342(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_343_555 <= heap_bh30_w127_8 & heap_bh30_w127_7 & heap_bh30_w127_6;
   CompressorIn_bh30_343_556 <= heap_bh30_w128_8 & heap_bh30_w128_7;
      Compressor_bh30_343: Compressor_23_3
      port map ( R => CompressorOut_bh30_343_343,
                 X0 => CompressorIn_bh30_343_555,
                 X1 => CompressorIn_bh30_343_556);
   heap_bh30_w127_10 <= CompressorOut_bh30_343_343(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w128_9 <= CompressorOut_bh30_343_343(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w129_9 <= CompressorOut_bh30_343_343(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_344_557 <= heap_bh30_w131_7 & heap_bh30_w131_6 & heap_bh30_w131_5;
   CompressorIn_bh30_344_558 <= heap_bh30_w132_6 & heap_bh30_w132_5;
      Compressor_bh30_344: Compressor_23_3
      port map ( R => CompressorOut_bh30_344_344,
                 X0 => CompressorIn_bh30_344_557,
                 X1 => CompressorIn_bh30_344_558);
   heap_bh30_w131_9 <= CompressorOut_bh30_344_344(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w132_7 <= CompressorOut_bh30_344_344(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w133_7 <= CompressorOut_bh30_344_344(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_345_559 <= heap_bh30_w133_6 & heap_bh30_w133_5 & heap_bh30_w133_4;
   CompressorIn_bh30_345_560 <= heap_bh30_w134_5 & heap_bh30_w134_4;
      Compressor_bh30_345: Compressor_23_3
      port map ( R => CompressorOut_bh30_345_345,
                 X0 => CompressorIn_bh30_345_559,
                 X1 => CompressorIn_bh30_345_560);
   heap_bh30_w133_8 <= CompressorOut_bh30_345_345(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w134_6 <= CompressorOut_bh30_345_345(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w135_7 <= CompressorOut_bh30_345_345(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_346_561 <= heap_bh30_w135_6 & heap_bh30_w135_5 & heap_bh30_w135_4;
   CompressorIn_bh30_346_562 <= heap_bh30_w136_5 & heap_bh30_w136_4;
      Compressor_bh30_346: Compressor_23_3
      port map ( R => CompressorOut_bh30_346_346,
                 X0 => CompressorIn_bh30_346_561,
                 X1 => CompressorIn_bh30_346_562);
   heap_bh30_w135_8 <= CompressorOut_bh30_346_346(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w136_6 <= CompressorOut_bh30_346_346(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w137_7 <= CompressorOut_bh30_346_346(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_347_563 <= heap_bh30_w137_6 & heap_bh30_w137_5 & heap_bh30_w137_4;
   CompressorIn_bh30_347_564 <= heap_bh30_w138_5 & heap_bh30_w138_4;
      Compressor_bh30_347: Compressor_23_3
      port map ( R => CompressorOut_bh30_347_347,
                 X0 => CompressorIn_bh30_347_563,
                 X1 => CompressorIn_bh30_347_564);
   heap_bh30_w137_8 <= CompressorOut_bh30_347_347(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w138_6 <= CompressorOut_bh30_347_347(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w139_7 <= CompressorOut_bh30_347_347(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_348_565 <= heap_bh30_w139_6 & heap_bh30_w139_5 & heap_bh30_w139_4;
   CompressorIn_bh30_348_566 <= heap_bh30_w140_5 & heap_bh30_w140_4;
      Compressor_bh30_348: Compressor_23_3
      port map ( R => CompressorOut_bh30_348_348,
                 X0 => CompressorIn_bh30_348_565,
                 X1 => CompressorIn_bh30_348_566);
   heap_bh30_w139_8 <= CompressorOut_bh30_348_348(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w140_6 <= CompressorOut_bh30_348_348(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w141_7 <= CompressorOut_bh30_348_348(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_349_567 <= heap_bh30_w141_6 & heap_bh30_w141_5 & heap_bh30_w141_4;
   CompressorIn_bh30_349_568 <= heap_bh30_w142_5 & heap_bh30_w142_4;
      Compressor_bh30_349: Compressor_23_3
      port map ( R => CompressorOut_bh30_349_349,
                 X0 => CompressorIn_bh30_349_567,
                 X1 => CompressorIn_bh30_349_568);
   heap_bh30_w141_8 <= CompressorOut_bh30_349_349(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w142_6 <= CompressorOut_bh30_349_349(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w143_7 <= CompressorOut_bh30_349_349(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_350_569 <= heap_bh30_w143_6 & heap_bh30_w143_5 & heap_bh30_w143_4;
   CompressorIn_bh30_350_570 <= heap_bh30_w144_5 & heap_bh30_w144_4;
      Compressor_bh30_350: Compressor_23_3
      port map ( R => CompressorOut_bh30_350_350,
                 X0 => CompressorIn_bh30_350_569,
                 X1 => CompressorIn_bh30_350_570);
   heap_bh30_w143_8 <= CompressorOut_bh30_350_350(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w144_6 <= CompressorOut_bh30_350_350(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w145_7 <= CompressorOut_bh30_350_350(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_351_571 <= heap_bh30_w145_6 & heap_bh30_w145_5 & heap_bh30_w145_4;
   CompressorIn_bh30_351_572 <= heap_bh30_w146_1 & heap_bh30_w146_0;
      Compressor_bh30_351: Compressor_23_3
      port map ( R => CompressorOut_bh30_351_351,
                 X0 => CompressorIn_bh30_351_571,
                 X1 => CompressorIn_bh30_351_572);
   heap_bh30_w145_8 <= CompressorOut_bh30_351_351(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w146_4 <= CompressorOut_bh30_351_351(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w147_5 <= CompressorOut_bh30_351_351(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_352_573 <= heap_bh30_w157_1 & heap_bh30_w157_0 & heap_bh30_w157_2;
   CompressorIn_bh30_352_574 <= heap_bh30_w158_1 & heap_bh30_w158_0;
      Compressor_bh30_352: Compressor_23_3
      port map ( R => CompressorOut_bh30_352_352,
                 X0 => CompressorIn_bh30_352_573,
                 X1 => CompressorIn_bh30_352_574);
   heap_bh30_w157_3 <= CompressorOut_bh30_352_352(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w158_2 <= CompressorOut_bh30_352_352(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w159_2 <= CompressorOut_bh30_352_352(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_353_575 <= heap_bh30_w14_7 & heap_bh30_w14_3 & heap_bh30_w14_8;
   CompressorIn_bh30_353_576(0) <= heap_bh30_w15_9;
      Compressor_bh30_353: Compressor_13_3
      port map ( R => CompressorOut_bh30_353_353,
                 X0 => CompressorIn_bh30_353_575,
                 X1 => CompressorIn_bh30_353_576);
   heap_bh30_w14_9 <= CompressorOut_bh30_353_353(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w15_10 <= CompressorOut_bh30_353_353(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w16_11 <= CompressorOut_bh30_353_353(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_354_577 <= heap_bh30_w36_14 & heap_bh30_w36_13 & heap_bh30_w36_12;
      Compressor_bh30_354: Compressor_3_2
      port map ( R => CompressorOut_bh30_354_354,
                 X0 => CompressorIn_bh30_354_577);
   heap_bh30_w36_16 <= CompressorOut_bh30_354_354(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w37_16 <= CompressorOut_bh30_354_354(1); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_355_578 <= heap_bh30_w39_14 & heap_bh30_w39_13 & heap_bh30_w39_12;
      Compressor_bh30_355: Compressor_3_2
      port map ( R => CompressorOut_bh30_355_355,
                 X0 => CompressorIn_bh30_355_578);
   heap_bh30_w39_16 <= CompressorOut_bh30_355_355(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w40_16 <= CompressorOut_bh30_355_355(1); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_356_579 <= heap_bh30_w42_14 & heap_bh30_w42_13 & heap_bh30_w42_12;
      Compressor_bh30_356: Compressor_3_2
      port map ( R => CompressorOut_bh30_356_356,
                 X0 => CompressorIn_bh30_356_579);
   heap_bh30_w42_16 <= CompressorOut_bh30_356_356(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w43_16 <= CompressorOut_bh30_356_356(1); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_357_580 <= heap_bh30_w47_14 & heap_bh30_w47_13 & heap_bh30_w47_12;
      Compressor_bh30_357: Compressor_3_2
      port map ( R => CompressorOut_bh30_357_357,
                 X0 => CompressorIn_bh30_357_580);
   heap_bh30_w47_16 <= CompressorOut_bh30_357_357(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w48_17 <= CompressorOut_bh30_357_357(1); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_358_581 <= heap_bh30_w52_16 & heap_bh30_w52_15 & heap_bh30_w52_14;
      Compressor_bh30_358: Compressor_3_2
      port map ( R => CompressorOut_bh30_358_358,
                 X0 => CompressorIn_bh30_358_581);
   heap_bh30_w52_19 <= CompressorOut_bh30_358_358(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w53_18 <= CompressorOut_bh30_358_358(1); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_359_582 <= heap_bh30_w55_16 & heap_bh30_w55_15 & heap_bh30_w55_14;
      Compressor_bh30_359: Compressor_3_2
      port map ( R => CompressorOut_bh30_359_359,
                 X0 => CompressorIn_bh30_359_582);
   heap_bh30_w55_19 <= CompressorOut_bh30_359_359(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w56_18 <= CompressorOut_bh30_359_359(1); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_360_583 <= heap_bh30_w58_16 & heap_bh30_w58_15 & heap_bh30_w58_14;
      Compressor_bh30_360: Compressor_3_2
      port map ( R => CompressorOut_bh30_360_360,
                 X0 => CompressorIn_bh30_360_583);
   heap_bh30_w58_19 <= CompressorOut_bh30_360_360(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w59_18 <= CompressorOut_bh30_360_360(1); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_361_584 <= heap_bh30_w61_16 & heap_bh30_w61_15 & heap_bh30_w61_14;
      Compressor_bh30_361: Compressor_3_2
      port map ( R => CompressorOut_bh30_361_361,
                 X0 => CompressorIn_bh30_361_584);
   heap_bh30_w61_19 <= CompressorOut_bh30_361_361(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w62_18 <= CompressorOut_bh30_361_361(1); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_362_585 <= heap_bh30_w64_16 & heap_bh30_w64_15 & heap_bh30_w64_14;
      Compressor_bh30_362: Compressor_3_2
      port map ( R => CompressorOut_bh30_362_362,
                 X0 => CompressorIn_bh30_362_585);
   heap_bh30_w64_19 <= CompressorOut_bh30_362_362(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w65_18 <= CompressorOut_bh30_362_362(1); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_363_586 <= heap_bh30_w69_17 & heap_bh30_w69_16 & heap_bh30_w69_15;
      Compressor_bh30_363: Compressor_3_2
      port map ( R => CompressorOut_bh30_363_363,
                 X0 => CompressorIn_bh30_363_586);
   heap_bh30_w69_21 <= CompressorOut_bh30_363_363(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w70_21 <= CompressorOut_bh30_363_363(1); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_364_587 <= heap_bh30_w108_9 & heap_bh30_w108_8 & heap_bh30_w108_7;
      Compressor_bh30_364: Compressor_3_2
      port map ( R => CompressorOut_bh30_364_364,
                 X0 => CompressorIn_bh30_364_587);
   heap_bh30_w108_12 <= CompressorOut_bh30_364_364(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w109_12 <= CompressorOut_bh30_364_364(1); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_365_588 <= heap_bh30_w110_9 & heap_bh30_w110_8 & heap_bh30_w110_7;
      Compressor_bh30_365: Compressor_3_2
      port map ( R => CompressorOut_bh30_365_365,
                 X0 => CompressorIn_bh30_365_588);
   heap_bh30_w110_11 <= CompressorOut_bh30_365_365(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w111_12 <= CompressorOut_bh30_365_365(1); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_366_589 <= heap_bh30_w74_15 & heap_bh30_w74_22 & heap_bh30_w74_21 & heap_bh30_w74_20;
   CompressorIn_bh30_366_590(0) <= heap_bh30_w75_23;
      Compressor_bh30_366: Compressor_14_3
      port map ( R => CompressorOut_bh30_366_366,
                 X0 => CompressorIn_bh30_366_589,
                 X1 => CompressorIn_bh30_366_590);
   heap_bh30_w74_23 <= CompressorOut_bh30_366_366(0); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w75_24 <= CompressorOut_bh30_366_366(1); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w76_23 <= CompressorOut_bh30_366_366(2); -- cycle= 0 cp= 3.97916e-09

   CompressorIn_bh30_367_591 <= heap_bh30_w77_15 & heap_bh30_w77_22 & heap_bh30_w77_21 & heap_bh30_w77_20;
   CompressorIn_bh30_367_592(0) <= heap_bh30_w78_23;
      Compressor_bh30_367: Compressor_14_3
      port map ( R => CompressorOut_bh30_367_367,
                 X0 => CompressorIn_bh30_367_591,
                 X1 => CompressorIn_bh30_367_592);
   heap_bh30_w77_23 <= CompressorOut_bh30_367_367(0); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w78_24 <= CompressorOut_bh30_367_367(1); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w79_23 <= CompressorOut_bh30_367_367(2); -- cycle= 0 cp= 3.97916e-09

   CompressorIn_bh30_368_593 <= heap_bh30_w80_15 & heap_bh30_w80_22 & heap_bh30_w80_21 & heap_bh30_w80_20;
   CompressorIn_bh30_368_594(0) <= heap_bh30_w81_23;
      Compressor_bh30_368: Compressor_14_3
      port map ( R => CompressorOut_bh30_368_368,
                 X0 => CompressorIn_bh30_368_593,
                 X1 => CompressorIn_bh30_368_594);
   heap_bh30_w80_23 <= CompressorOut_bh30_368_368(0); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w81_24 <= CompressorOut_bh30_368_368(1); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w82_23 <= CompressorOut_bh30_368_368(2); -- cycle= 0 cp= 3.97916e-09

   CompressorIn_bh30_369_595 <= heap_bh30_w83_15 & heap_bh30_w83_22 & heap_bh30_w83_21 & heap_bh30_w83_20;
   CompressorIn_bh30_369_596(0) <= heap_bh30_w84_23;
      Compressor_bh30_369: Compressor_14_3
      port map ( R => CompressorOut_bh30_369_369,
                 X0 => CompressorIn_bh30_369_595,
                 X1 => CompressorIn_bh30_369_596);
   heap_bh30_w83_23 <= CompressorOut_bh30_369_369(0); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w84_24 <= CompressorOut_bh30_369_369(1); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w85_23 <= CompressorOut_bh30_369_369(2); -- cycle= 0 cp= 3.97916e-09

   CompressorIn_bh30_370_597 <= heap_bh30_w86_15 & heap_bh30_w86_22 & heap_bh30_w86_21 & heap_bh30_w86_20;
   CompressorIn_bh30_370_598(0) <= heap_bh30_w87_23;
      Compressor_bh30_370: Compressor_14_3
      port map ( R => CompressorOut_bh30_370_370,
                 X0 => CompressorIn_bh30_370_597,
                 X1 => CompressorIn_bh30_370_598);
   heap_bh30_w86_23 <= CompressorOut_bh30_370_370(0); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w87_24 <= CompressorOut_bh30_370_370(1); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w88_23 <= CompressorOut_bh30_370_370(2); -- cycle= 0 cp= 3.97916e-09

   CompressorIn_bh30_371_599 <= heap_bh30_w89_15 & heap_bh30_w89_22 & heap_bh30_w89_21 & heap_bh30_w89_20;
   CompressorIn_bh30_371_600(0) <= heap_bh30_w90_22;
      Compressor_bh30_371: Compressor_14_3
      port map ( R => CompressorOut_bh30_371_371,
                 X0 => CompressorIn_bh30_371_599,
                 X1 => CompressorIn_bh30_371_600);
   heap_bh30_w89_23 <= CompressorOut_bh30_371_371(0); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w90_23 <= CompressorOut_bh30_371_371(1); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w91_21 <= CompressorOut_bh30_371_371(2); -- cycle= 0 cp= 3.97916e-09

   CompressorIn_bh30_372_601 <= heap_bh30_w92_11 & heap_bh30_w92_18 & heap_bh30_w92_17 & heap_bh30_w92_16;
   CompressorIn_bh30_372_602(0) <= heap_bh30_w93_17;
      Compressor_bh30_372: Compressor_14_3
      port map ( R => CompressorOut_bh30_372_372,
                 X0 => CompressorIn_bh30_372_601,
                 X1 => CompressorIn_bh30_372_602);
   heap_bh30_w92_19 <= CompressorOut_bh30_372_372(0); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w93_18 <= CompressorOut_bh30_372_372(1); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w94_16 <= CompressorOut_bh30_372_372(2); -- cycle= 0 cp= 3.97916e-09

   CompressorIn_bh30_373_603 <= heap_bh30_w96_8 & heap_bh30_w96_13 & heap_bh30_w96_12 & heap_bh30_w96_11;
   CompressorIn_bh30_373_604(0) <= heap_bh30_w97_13;
      Compressor_bh30_373: Compressor_14_3
      port map ( R => CompressorOut_bh30_373_373,
                 X0 => CompressorIn_bh30_373_603,
                 X1 => CompressorIn_bh30_373_604);
   heap_bh30_w96_14 <= CompressorOut_bh30_373_373(0); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w97_14 <= CompressorOut_bh30_373_373(1); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w98_14 <= CompressorOut_bh30_373_373(2); -- cycle= 0 cp= 3.97916e-09

   CompressorIn_bh30_374_605 <= heap_bh30_w10_8 & heap_bh30_w10_4 & heap_bh30_w10_9;
   CompressorIn_bh30_374_606 <= heap_bh30_w11_7 & heap_bh30_w11_3;
      Compressor_bh30_374: Compressor_23_3
      port map ( R => CompressorOut_bh30_374_374,
                 X0 => CompressorIn_bh30_374_605,
                 X1 => CompressorIn_bh30_374_606);
   heap_bh30_w10_10 <= CompressorOut_bh30_374_374(0); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w11_8 <= CompressorOut_bh30_374_374(1); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w12_10 <= CompressorOut_bh30_374_374(2); -- cycle= 0 cp= 3.97916e-09

   CompressorIn_bh30_375_607 <= heap_bh30_w16_4 & heap_bh30_w16_10 & heap_bh30_w16_11;
   CompressorIn_bh30_375_608 <= heap_bh30_w17_10 & heap_bh30_w17_9;
      Compressor_bh30_375: Compressor_23_3
      port map ( R => CompressorOut_bh30_375_375,
                 X0 => CompressorIn_bh30_375_607,
                 X1 => CompressorIn_bh30_375_608);
   heap_bh30_w16_12 <= CompressorOut_bh30_375_375(0); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w17_11 <= CompressorOut_bh30_375_375(1); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w18_12 <= CompressorOut_bh30_375_375(2); -- cycle= 0 cp= 3.97916e-09

   CompressorIn_bh30_376_609 <= heap_bh30_w35_12 & heap_bh30_w35_11 & heap_bh30_w35_14;
   CompressorIn_bh30_376_610 <= heap_bh30_w36_16 & heap_bh30_w36_15;
      Compressor_bh30_376: Compressor_23_3
      port map ( R => CompressorOut_bh30_376_376,
                 X0 => CompressorIn_bh30_376_609,
                 X1 => CompressorIn_bh30_376_610);
   heap_bh30_w35_15 <= CompressorOut_bh30_376_376(0); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w36_17 <= CompressorOut_bh30_376_376(1); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w37_17 <= CompressorOut_bh30_376_376(2); -- cycle= 0 cp= 3.97916e-09

   CompressorIn_bh30_377_611 <= heap_bh30_w38_12 & heap_bh30_w38_11 & heap_bh30_w38_14;
   CompressorIn_bh30_377_612 <= heap_bh30_w39_16 & heap_bh30_w39_15;
      Compressor_bh30_377: Compressor_23_3
      port map ( R => CompressorOut_bh30_377_377,
                 X0 => CompressorIn_bh30_377_611,
                 X1 => CompressorIn_bh30_377_612);
   heap_bh30_w38_15 <= CompressorOut_bh30_377_377(0); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w39_17 <= CompressorOut_bh30_377_377(1); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w40_17 <= CompressorOut_bh30_377_377(2); -- cycle= 0 cp= 3.97916e-09

   CompressorIn_bh30_378_613 <= heap_bh30_w41_12 & heap_bh30_w41_11 & heap_bh30_w41_14;
   CompressorIn_bh30_378_614 <= heap_bh30_w42_16 & heap_bh30_w42_15;
      Compressor_bh30_378: Compressor_23_3
      port map ( R => CompressorOut_bh30_378_378,
                 X0 => CompressorIn_bh30_378_613,
                 X1 => CompressorIn_bh30_378_614);
   heap_bh30_w41_15 <= CompressorOut_bh30_378_378(0); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w42_17 <= CompressorOut_bh30_378_378(1); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w43_17 <= CompressorOut_bh30_378_378(2); -- cycle= 0 cp= 3.97916e-09

   CompressorIn_bh30_379_615 <= heap_bh30_w44_12 & heap_bh30_w44_11 & heap_bh30_w44_14;
   CompressorIn_bh30_379_616 <= heap_bh30_w45_16 & heap_bh30_w45_15;
      Compressor_bh30_379: Compressor_23_3
      port map ( R => CompressorOut_bh30_379_379,
                 X0 => CompressorIn_bh30_379_615,
                 X1 => CompressorIn_bh30_379_616);
   heap_bh30_w44_15 <= CompressorOut_bh30_379_379(0); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w45_17 <= CompressorOut_bh30_379_379(1); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w46_16 <= CompressorOut_bh30_379_379(2); -- cycle= 0 cp= 3.97916e-09

   CompressorIn_bh30_380_617 <= heap_bh30_w49_14 & heap_bh30_w49_13 & heap_bh30_w49_16;
   CompressorIn_bh30_380_618 <= heap_bh30_w50_17 & heap_bh30_w50_16;
      Compressor_bh30_380: Compressor_23_3
      port map ( R => CompressorOut_bh30_380_380,
                 X0 => CompressorIn_bh30_380_617,
                 X1 => CompressorIn_bh30_380_618);
   heap_bh30_w49_17 <= CompressorOut_bh30_380_380(0); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w50_18 <= CompressorOut_bh30_380_380(1); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w51_19 <= CompressorOut_bh30_380_380(2); -- cycle= 0 cp= 3.97916e-09

   CompressorIn_bh30_381_619 <= heap_bh30_w52_19 & heap_bh30_w52_18 & heap_bh30_w52_17;
   CompressorIn_bh30_381_620 <= heap_bh30_w53_18 & heap_bh30_w53_17;
      Compressor_bh30_381: Compressor_23_3
      port map ( R => CompressorOut_bh30_381_381,
                 X0 => CompressorIn_bh30_381_619,
                 X1 => CompressorIn_bh30_381_620);
   heap_bh30_w52_20 <= CompressorOut_bh30_381_381(0); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w53_19 <= CompressorOut_bh30_381_381(1); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w54_19 <= CompressorOut_bh30_381_381(2); -- cycle= 0 cp= 3.97916e-09

   CompressorIn_bh30_382_621 <= heap_bh30_w55_19 & heap_bh30_w55_18 & heap_bh30_w55_17;
   CompressorIn_bh30_382_622 <= heap_bh30_w56_18 & heap_bh30_w56_17;
      Compressor_bh30_382: Compressor_23_3
      port map ( R => CompressorOut_bh30_382_382,
                 X0 => CompressorIn_bh30_382_621,
                 X1 => CompressorIn_bh30_382_622);
   heap_bh30_w55_20 <= CompressorOut_bh30_382_382(0); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w56_19 <= CompressorOut_bh30_382_382(1); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w57_19 <= CompressorOut_bh30_382_382(2); -- cycle= 0 cp= 3.97916e-09

   CompressorIn_bh30_383_623 <= heap_bh30_w58_19 & heap_bh30_w58_18 & heap_bh30_w58_17;
   CompressorIn_bh30_383_624 <= heap_bh30_w59_18 & heap_bh30_w59_17;
      Compressor_bh30_383: Compressor_23_3
      port map ( R => CompressorOut_bh30_383_383,
                 X0 => CompressorIn_bh30_383_623,
                 X1 => CompressorIn_bh30_383_624);
   heap_bh30_w58_20 <= CompressorOut_bh30_383_383(0); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w59_19 <= CompressorOut_bh30_383_383(1); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w60_19 <= CompressorOut_bh30_383_383(2); -- cycle= 0 cp= 3.97916e-09

   CompressorIn_bh30_384_625 <= heap_bh30_w61_19 & heap_bh30_w61_18 & heap_bh30_w61_17;
   CompressorIn_bh30_384_626 <= heap_bh30_w62_18 & heap_bh30_w62_17;
      Compressor_bh30_384: Compressor_23_3
      port map ( R => CompressorOut_bh30_384_384,
                 X0 => CompressorIn_bh30_384_625,
                 X1 => CompressorIn_bh30_384_626);
   heap_bh30_w61_20 <= CompressorOut_bh30_384_384(0); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w62_19 <= CompressorOut_bh30_384_384(1); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w63_19 <= CompressorOut_bh30_384_384(2); -- cycle= 0 cp= 3.97916e-09

   CompressorIn_bh30_385_627 <= heap_bh30_w64_19 & heap_bh30_w64_18 & heap_bh30_w64_17;
   CompressorIn_bh30_385_628 <= heap_bh30_w65_18 & heap_bh30_w65_17;
      Compressor_bh30_385: Compressor_23_3
      port map ( R => CompressorOut_bh30_385_385,
                 X0 => CompressorIn_bh30_385_627,
                 X1 => CompressorIn_bh30_385_628);
   heap_bh30_w64_20 <= CompressorOut_bh30_385_385(0); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w65_19 <= CompressorOut_bh30_385_385(1); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w66_19 <= CompressorOut_bh30_385_385(2); -- cycle= 0 cp= 3.97916e-09

   CompressorIn_bh30_386_629 <= heap_bh30_w67_20 & heap_bh30_w67_19 & heap_bh30_w67_18;
   CompressorIn_bh30_386_630 <= heap_bh30_w68_19 & heap_bh30_w68_18;
      Compressor_bh30_386: Compressor_23_3
      port map ( R => CompressorOut_bh30_386_386,
                 X0 => CompressorIn_bh30_386_629,
                 X1 => CompressorIn_bh30_386_630);
   heap_bh30_w67_21 <= CompressorOut_bh30_386_386(0); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w68_20 <= CompressorOut_bh30_386_386(1); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w69_22 <= CompressorOut_bh30_386_386(2); -- cycle= 0 cp= 3.97916e-09

   CompressorIn_bh30_387_631 <= heap_bh30_w69_21 & heap_bh30_w69_20 & heap_bh30_w69_19;
   CompressorIn_bh30_387_632 <= heap_bh30_w70_21 & heap_bh30_w70_20;
      Compressor_bh30_387: Compressor_23_3
      port map ( R => CompressorOut_bh30_387_387,
                 X0 => CompressorIn_bh30_387_631,
                 X1 => CompressorIn_bh30_387_632);
   heap_bh30_w69_23 <= CompressorOut_bh30_387_387(0); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w70_22 <= CompressorOut_bh30_387_387(1); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w71_22 <= CompressorOut_bh30_387_387(2); -- cycle= 0 cp= 3.97916e-09

   CompressorIn_bh30_388_633 <= heap_bh30_w72_23 & heap_bh30_w72_22 & heap_bh30_w72_21;
   CompressorIn_bh30_388_634 <= heap_bh30_w73_22 & heap_bh30_w73_21;
      Compressor_bh30_388: Compressor_23_3
      port map ( R => CompressorOut_bh30_388_388,
                 X0 => CompressorIn_bh30_388_633,
                 X1 => CompressorIn_bh30_388_634);
   heap_bh30_w72_24 <= CompressorOut_bh30_388_388(0); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w73_23 <= CompressorOut_bh30_388_388(1); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w74_24 <= CompressorOut_bh30_388_388(2); -- cycle= 0 cp= 3.97916e-09

   CompressorIn_bh30_389_635 <= heap_bh30_w94_15 & heap_bh30_w94_14 & heap_bh30_w94_13;
   CompressorIn_bh30_389_636 <= heap_bh30_w95_14 & heap_bh30_w95_13;
      Compressor_bh30_389: Compressor_23_3
      port map ( R => CompressorOut_bh30_389_389,
                 X0 => CompressorIn_bh30_389_635,
                 X1 => CompressorIn_bh30_389_636);
   heap_bh30_w94_17 <= CompressorOut_bh30_389_389(0); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w95_15 <= CompressorOut_bh30_389_389(1); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w96_15 <= CompressorOut_bh30_389_389(2); -- cycle= 0 cp= 3.97916e-09

   CompressorIn_bh30_390_637 <= heap_bh30_w98_13 & heap_bh30_w98_12 & heap_bh30_w98_11;
   CompressorIn_bh30_390_638 <= heap_bh30_w99_13 & heap_bh30_w99_12;
      Compressor_bh30_390: Compressor_23_3
      port map ( R => CompressorOut_bh30_390_390,
                 X0 => CompressorIn_bh30_390_637,
                 X1 => CompressorIn_bh30_390_638);
   heap_bh30_w98_15 <= CompressorOut_bh30_390_390(0); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w99_14 <= CompressorOut_bh30_390_390(1); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w100_14 <= CompressorOut_bh30_390_390(2); -- cycle= 0 cp= 3.97916e-09

   CompressorIn_bh30_391_639 <= heap_bh30_w100_13 & heap_bh30_w100_12 & heap_bh30_w100_11;
   CompressorIn_bh30_391_640 <= heap_bh30_w101_13 & heap_bh30_w101_12;
      Compressor_bh30_391: Compressor_23_3
      port map ( R => CompressorOut_bh30_391_391,
                 X0 => CompressorIn_bh30_391_639,
                 X1 => CompressorIn_bh30_391_640);
   heap_bh30_w100_15 <= CompressorOut_bh30_391_391(0); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w101_14 <= CompressorOut_bh30_391_391(1); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w102_14 <= CompressorOut_bh30_391_391(2); -- cycle= 0 cp= 3.97916e-09

   CompressorIn_bh30_392_641 <= heap_bh30_w102_13 & heap_bh30_w102_12 & heap_bh30_w102_11;
   CompressorIn_bh30_392_642 <= heap_bh30_w103_13 & heap_bh30_w103_12;
      Compressor_bh30_392: Compressor_23_3
      port map ( R => CompressorOut_bh30_392_392,
                 X0 => CompressorIn_bh30_392_641,
                 X1 => CompressorIn_bh30_392_642);
   heap_bh30_w102_15 <= CompressorOut_bh30_392_392(0); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w103_14 <= CompressorOut_bh30_392_392(1); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w104_14 <= CompressorOut_bh30_392_392(2); -- cycle= 0 cp= 3.97916e-09

   CompressorIn_bh30_393_643 <= heap_bh30_w104_13 & heap_bh30_w104_12 & heap_bh30_w104_11;
   CompressorIn_bh30_393_644 <= heap_bh30_w105_13 & heap_bh30_w105_12;
      Compressor_bh30_393: Compressor_23_3
      port map ( R => CompressorOut_bh30_393_393,
                 X0 => CompressorIn_bh30_393_643,
                 X1 => CompressorIn_bh30_393_644);
   heap_bh30_w104_15 <= CompressorOut_bh30_393_393(0); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w105_14 <= CompressorOut_bh30_393_393(1); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w106_14 <= CompressorOut_bh30_393_393(2); -- cycle= 0 cp= 3.97916e-09

   CompressorIn_bh30_394_645 <= heap_bh30_w106_13 & heap_bh30_w106_12 & heap_bh30_w106_11;
   CompressorIn_bh30_394_646 <= heap_bh30_w107_13 & heap_bh30_w107_12;
      Compressor_bh30_394: Compressor_23_3
      port map ( R => CompressorOut_bh30_394_394,
                 X0 => CompressorIn_bh30_394_645,
                 X1 => CompressorIn_bh30_394_646);
   heap_bh30_w106_15 <= CompressorOut_bh30_394_394(0); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w107_14 <= CompressorOut_bh30_394_394(1); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w108_13 <= CompressorOut_bh30_394_394(2); -- cycle= 0 cp= 3.97916e-09

   CompressorIn_bh30_395_647 <= heap_bh30_w108_12 & heap_bh30_w108_11 & heap_bh30_w108_10;
   CompressorIn_bh30_395_648 <= heap_bh30_w109_12 & heap_bh30_w109_11;
      Compressor_bh30_395: Compressor_23_3
      port map ( R => CompressorOut_bh30_395_395,
                 X0 => CompressorIn_bh30_395_647,
                 X1 => CompressorIn_bh30_395_648);
   heap_bh30_w108_14 <= CompressorOut_bh30_395_395(0); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w109_13 <= CompressorOut_bh30_395_395(1); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w110_12 <= CompressorOut_bh30_395_395(2); -- cycle= 0 cp= 3.97916e-09

   CompressorIn_bh30_396_649 <= heap_bh30_w111_12 & heap_bh30_w111_11 & heap_bh30_w111_10;
   CompressorIn_bh30_396_650 <= heap_bh30_w112_7 & heap_bh30_w112_6;
      Compressor_bh30_396: Compressor_23_3
      port map ( R => CompressorOut_bh30_396_396,
                 X0 => CompressorIn_bh30_396_649,
                 X1 => CompressorIn_bh30_396_650);
   heap_bh30_w111_13 <= CompressorOut_bh30_396_396(0); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w112_10 <= CompressorOut_bh30_396_396(1); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w113_11 <= CompressorOut_bh30_396_396(2); -- cycle= 0 cp= 3.97916e-09

   CompressorIn_bh30_397_651 <= heap_bh30_w130_6 & heap_bh30_w130_5 & heap_bh30_w130_8;
   CompressorIn_bh30_397_652 <= heap_bh30_w131_9 & heap_bh30_w131_8;
      Compressor_bh30_397: Compressor_23_3
      port map ( R => CompressorOut_bh30_397_397,
                 X0 => CompressorIn_bh30_397_651,
                 X1 => CompressorIn_bh30_397_652);
   heap_bh30_w130_9 <= CompressorOut_bh30_397_397(0); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w131_10 <= CompressorOut_bh30_397_397(1); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w132_8 <= CompressorOut_bh30_397_397(2); -- cycle= 0 cp= 3.97916e-09

   CompressorIn_bh30_398_653 <= heap_bh30_w147_4 & heap_bh30_w147_3 & heap_bh30_w147_5;
   CompressorIn_bh30_398_654 <= heap_bh30_w148_0 & heap_bh30_w148_3;
      Compressor_bh30_398: Compressor_23_3
      port map ( R => CompressorOut_bh30_398_398,
                 X0 => CompressorIn_bh30_398_653,
                 X1 => CompressorIn_bh30_398_654);
   heap_bh30_w147_6 <= CompressorOut_bh30_398_398(0); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w148_4 <= CompressorOut_bh30_398_398(1); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w149_5 <= CompressorOut_bh30_398_398(2); -- cycle= 0 cp= 3.97916e-09

   CompressorIn_bh30_399_655 <= heap_bh30_w159_1 & heap_bh30_w159_0 & heap_bh30_w159_2;
   CompressorIn_bh30_399_656 <= heap_bh30_w160_1 & heap_bh30_w160_0;
      Compressor_bh30_399: Compressor_23_3
      port map ( R => CompressorOut_bh30_399_399,
                 X0 => CompressorIn_bh30_399_655,
                 X1 => CompressorIn_bh30_399_656);
   heap_bh30_w159_3 <= CompressorOut_bh30_399_399(0); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w160_2 <= CompressorOut_bh30_399_399(1); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w161_2 <= CompressorOut_bh30_399_399(2); -- cycle= 0 cp= 3.97916e-09

   CompressorIn_bh30_400_657 <= heap_bh30_w21_11 & heap_bh30_w21_10 & heap_bh30_w21_12;
   CompressorIn_bh30_400_658(0) <= heap_bh30_w22_11;
      Compressor_bh30_400: Compressor_13_3
      port map ( R => CompressorOut_bh30_400_400,
                 X0 => CompressorIn_bh30_400_657,
                 X1 => CompressorIn_bh30_400_658);
   heap_bh30_w21_13 <= CompressorOut_bh30_400_400(0); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w22_12 <= CompressorOut_bh30_400_400(1); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w23_13 <= CompressorOut_bh30_400_400(2); -- cycle= 0 cp= 3.97916e-09

   CompressorIn_bh30_401_659 <= heap_bh30_w24_12 & heap_bh30_w24_11 & heap_bh30_w24_13;
   CompressorIn_bh30_401_660(0) <= heap_bh30_w25_14;
      Compressor_bh30_401: Compressor_13_3
      port map ( R => CompressorOut_bh30_401_401,
                 X0 => CompressorIn_bh30_401_659,
                 X1 => CompressorIn_bh30_401_660);
   heap_bh30_w24_14 <= CompressorOut_bh30_401_401(0); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w25_15 <= CompressorOut_bh30_401_401(1); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w26_14 <= CompressorOut_bh30_401_401(2); -- cycle= 0 cp= 3.97916e-09

   CompressorIn_bh30_402_661 <= heap_bh30_w27_12 & heap_bh30_w27_11 & heap_bh30_w27_13;
   CompressorIn_bh30_402_662(0) <= heap_bh30_w28_14;
      Compressor_bh30_402: Compressor_13_3
      port map ( R => CompressorOut_bh30_402_402,
                 X0 => CompressorIn_bh30_402_661,
                 X1 => CompressorIn_bh30_402_662);
   heap_bh30_w27_14 <= CompressorOut_bh30_402_402(0); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w28_15 <= CompressorOut_bh30_402_402(1); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w29_14 <= CompressorOut_bh30_402_402(2); -- cycle= 0 cp= 3.97916e-09

   CompressorIn_bh30_403_663 <= heap_bh30_w30_12 & heap_bh30_w30_11 & heap_bh30_w30_13;
   CompressorIn_bh30_403_664(0) <= heap_bh30_w31_14;
      Compressor_bh30_403: Compressor_13_3
      port map ( R => CompressorOut_bh30_403_403,
                 X0 => CompressorIn_bh30_403_663,
                 X1 => CompressorIn_bh30_403_664);
   heap_bh30_w30_14 <= CompressorOut_bh30_403_403(0); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w31_15 <= CompressorOut_bh30_403_403(1); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w32_14 <= CompressorOut_bh30_403_403(2); -- cycle= 0 cp= 3.97916e-09

   CompressorIn_bh30_404_665 <= heap_bh30_w33_13 & heap_bh30_w33_12 & heap_bh30_w33_14;
   CompressorIn_bh30_404_666(0) <= heap_bh30_w34_15;
      Compressor_bh30_404: Compressor_13_3
      port map ( R => CompressorOut_bh30_404_404,
                 X0 => CompressorIn_bh30_404_665,
                 X1 => CompressorIn_bh30_404_666);
   heap_bh30_w33_15 <= CompressorOut_bh30_404_404(0); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w34_16 <= CompressorOut_bh30_404_404(1); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w35_16 <= CompressorOut_bh30_404_404(2); -- cycle= 0 cp= 3.97916e-09

   CompressorIn_bh30_405_667 <= heap_bh30_w76_22 & heap_bh30_w76_21 & heap_bh30_w76_20;
      Compressor_bh30_405: Compressor_3_2
      port map ( R => CompressorOut_bh30_405_405,
                 X0 => CompressorIn_bh30_405_667);
   heap_bh30_w76_24 <= CompressorOut_bh30_405_405(0); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w77_24 <= CompressorOut_bh30_405_405(1); -- cycle= 0 cp= 3.97916e-09

   CompressorIn_bh30_406_668 <= heap_bh30_w79_22 & heap_bh30_w79_21 & heap_bh30_w79_20;
      Compressor_bh30_406: Compressor_3_2
      port map ( R => CompressorOut_bh30_406_406,
                 X0 => CompressorIn_bh30_406_668);
   heap_bh30_w79_24 <= CompressorOut_bh30_406_406(0); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w80_24 <= CompressorOut_bh30_406_406(1); -- cycle= 0 cp= 3.97916e-09

   CompressorIn_bh30_407_669 <= heap_bh30_w82_22 & heap_bh30_w82_21 & heap_bh30_w82_20;
      Compressor_bh30_407: Compressor_3_2
      port map ( R => CompressorOut_bh30_407_407,
                 X0 => CompressorIn_bh30_407_669);
   heap_bh30_w82_24 <= CompressorOut_bh30_407_407(0); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w83_24 <= CompressorOut_bh30_407_407(1); -- cycle= 0 cp= 3.97916e-09

   CompressorIn_bh30_408_670 <= heap_bh30_w85_22 & heap_bh30_w85_21 & heap_bh30_w85_20;
      Compressor_bh30_408: Compressor_3_2
      port map ( R => CompressorOut_bh30_408_408,
                 X0 => CompressorIn_bh30_408_670);
   heap_bh30_w85_24 <= CompressorOut_bh30_408_408(0); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w86_24 <= CompressorOut_bh30_408_408(1); -- cycle= 0 cp= 3.97916e-09

   CompressorIn_bh30_409_671 <= heap_bh30_w88_22 & heap_bh30_w88_21 & heap_bh30_w88_20;
      Compressor_bh30_409: Compressor_3_2
      port map ( R => CompressorOut_bh30_409_409,
                 X0 => CompressorIn_bh30_409_671);
   heap_bh30_w88_24 <= CompressorOut_bh30_409_409(0); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w89_24 <= CompressorOut_bh30_409_409(1); -- cycle= 0 cp= 3.97916e-09

   CompressorIn_bh30_410_672 <= heap_bh30_w91_20 & heap_bh30_w91_19 & heap_bh30_w91_18;
      Compressor_bh30_410: Compressor_3_2
      port map ( R => CompressorOut_bh30_410_410,
                 X0 => CompressorIn_bh30_410_672);
   heap_bh30_w91_22 <= CompressorOut_bh30_410_410(0); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w92_20 <= CompressorOut_bh30_410_410(1); -- cycle= 0 cp= 3.97916e-09

   CompressorIn_bh30_411_673 <= heap_bh30_w46_12 & heap_bh30_w46_15 & heap_bh30_w46_16;
   CompressorIn_bh30_411_674 <= heap_bh30_w47_16 & heap_bh30_w47_15;
      Compressor_bh30_411: Compressor_23_3
      port map ( R => CompressorOut_bh30_411_411,
                 X0 => CompressorIn_bh30_411_673,
                 X1 => CompressorIn_bh30_411_674);
   heap_bh30_w46_17 <= CompressorOut_bh30_411_411(0); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w47_17 <= CompressorOut_bh30_411_411(1); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w48_18 <= CompressorOut_bh30_411_411(2); -- cycle= 0 cp= 4.50988e-09

   CompressorIn_bh30_412_675 <= heap_bh30_w75_22 & heap_bh30_w75_21 & heap_bh30_w75_24;
   CompressorIn_bh30_412_676 <= heap_bh30_w76_24 & heap_bh30_w76_23;
      Compressor_bh30_412: Compressor_23_3
      port map ( R => CompressorOut_bh30_412_412,
                 X0 => CompressorIn_bh30_412_675,
                 X1 => CompressorIn_bh30_412_676);
   heap_bh30_w75_25 <= CompressorOut_bh30_412_412(0); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w76_25 <= CompressorOut_bh30_412_412(1); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w77_25 <= CompressorOut_bh30_412_412(2); -- cycle= 0 cp= 4.50988e-09

   CompressorIn_bh30_413_677 <= heap_bh30_w78_22 & heap_bh30_w78_21 & heap_bh30_w78_24;
   CompressorIn_bh30_413_678 <= heap_bh30_w79_24 & heap_bh30_w79_23;
      Compressor_bh30_413: Compressor_23_3
      port map ( R => CompressorOut_bh30_413_413,
                 X0 => CompressorIn_bh30_413_677,
                 X1 => CompressorIn_bh30_413_678);
   heap_bh30_w78_25 <= CompressorOut_bh30_413_413(0); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w79_25 <= CompressorOut_bh30_413_413(1); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w80_25 <= CompressorOut_bh30_413_413(2); -- cycle= 0 cp= 4.50988e-09

   CompressorIn_bh30_414_679 <= heap_bh30_w81_22 & heap_bh30_w81_21 & heap_bh30_w81_24;
   CompressorIn_bh30_414_680 <= heap_bh30_w82_24 & heap_bh30_w82_23;
      Compressor_bh30_414: Compressor_23_3
      port map ( R => CompressorOut_bh30_414_414,
                 X0 => CompressorIn_bh30_414_679,
                 X1 => CompressorIn_bh30_414_680);
   heap_bh30_w81_25 <= CompressorOut_bh30_414_414(0); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w82_25 <= CompressorOut_bh30_414_414(1); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w83_25 <= CompressorOut_bh30_414_414(2); -- cycle= 0 cp= 4.50988e-09

   CompressorIn_bh30_415_681 <= heap_bh30_w84_22 & heap_bh30_w84_21 & heap_bh30_w84_24;
   CompressorIn_bh30_415_682 <= heap_bh30_w85_24 & heap_bh30_w85_23;
      Compressor_bh30_415: Compressor_23_3
      port map ( R => CompressorOut_bh30_415_415,
                 X0 => CompressorIn_bh30_415_681,
                 X1 => CompressorIn_bh30_415_682);
   heap_bh30_w84_25 <= CompressorOut_bh30_415_415(0); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w85_25 <= CompressorOut_bh30_415_415(1); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w86_25 <= CompressorOut_bh30_415_415(2); -- cycle= 0 cp= 4.50988e-09

   CompressorIn_bh30_416_683 <= heap_bh30_w87_22 & heap_bh30_w87_21 & heap_bh30_w87_24;
   CompressorIn_bh30_416_684 <= heap_bh30_w88_24 & heap_bh30_w88_23;
      Compressor_bh30_416: Compressor_23_3
      port map ( R => CompressorOut_bh30_416_416,
                 X0 => CompressorIn_bh30_416_683,
                 X1 => CompressorIn_bh30_416_684);
   heap_bh30_w87_25 <= CompressorOut_bh30_416_416(0); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w88_25 <= CompressorOut_bh30_416_416(1); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w89_25 <= CompressorOut_bh30_416_416(2); -- cycle= 0 cp= 4.50988e-09

   CompressorIn_bh30_417_685 <= heap_bh30_w90_21 & heap_bh30_w90_20 & heap_bh30_w90_23;
   CompressorIn_bh30_417_686 <= heap_bh30_w91_22 & heap_bh30_w91_21;
      Compressor_bh30_417: Compressor_23_3
      port map ( R => CompressorOut_bh30_417_417,
                 X0 => CompressorIn_bh30_417_685,
                 X1 => CompressorIn_bh30_417_686);
   heap_bh30_w90_24 <= CompressorOut_bh30_417_417(0); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w91_23 <= CompressorOut_bh30_417_417(1); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w92_21 <= CompressorOut_bh30_417_417(2); -- cycle= 0 cp= 4.50988e-09

   CompressorIn_bh30_418_687 <= heap_bh30_w93_16 & heap_bh30_w93_15 & heap_bh30_w93_18;
   CompressorIn_bh30_418_688 <= heap_bh30_w94_17 & heap_bh30_w94_16;
      Compressor_bh30_418: Compressor_23_3
      port map ( R => CompressorOut_bh30_418_418,
                 X0 => CompressorIn_bh30_418_687,
                 X1 => CompressorIn_bh30_418_688);
   heap_bh30_w93_19 <= CompressorOut_bh30_418_418(0); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w94_18 <= CompressorOut_bh30_418_418(1); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w95_16 <= CompressorOut_bh30_418_418(2); -- cycle= 0 cp= 4.50988e-09

   CompressorIn_bh30_419_689 <= heap_bh30_w97_12 & heap_bh30_w97_11 & heap_bh30_w97_14;
   CompressorIn_bh30_419_690 <= heap_bh30_w98_15 & heap_bh30_w98_14;
      Compressor_bh30_419: Compressor_23_3
      port map ( R => CompressorOut_bh30_419_419,
                 X0 => CompressorIn_bh30_419_689,
                 X1 => CompressorIn_bh30_419_690);
   heap_bh30_w97_15 <= CompressorOut_bh30_419_419(0); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w98_16 <= CompressorOut_bh30_419_419(1); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w99_15 <= CompressorOut_bh30_419_419(2); -- cycle= 0 cp= 4.50988e-09

   CompressorIn_bh30_420_691 <= heap_bh30_w113_10 & heap_bh30_w113_9 & heap_bh30_w113_11;
   CompressorIn_bh30_420_692 <= heap_bh30_w114_6 & heap_bh30_w114_9;
      Compressor_bh30_420: Compressor_23_3
      port map ( R => CompressorOut_bh30_420_420,
                 X0 => CompressorIn_bh30_420_691,
                 X1 => CompressorIn_bh30_420_692);
   heap_bh30_w113_12 <= CompressorOut_bh30_420_420(0); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w114_10 <= CompressorOut_bh30_420_420(1); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w115_11 <= CompressorOut_bh30_420_420(2); -- cycle= 0 cp= 4.50988e-09

   CompressorIn_bh30_421_693 <= heap_bh30_w132_4 & heap_bh30_w132_7 & heap_bh30_w132_8;
   CompressorIn_bh30_421_694 <= heap_bh30_w133_8 & heap_bh30_w133_7;
      Compressor_bh30_421: Compressor_23_3
      port map ( R => CompressorOut_bh30_421_421,
                 X0 => CompressorIn_bh30_421_693,
                 X1 => CompressorIn_bh30_421_694);
   heap_bh30_w132_9 <= CompressorOut_bh30_421_421(0); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w133_9 <= CompressorOut_bh30_421_421(1); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w134_7 <= CompressorOut_bh30_421_421(2); -- cycle= 0 cp= 4.50988e-09

   CompressorIn_bh30_422_695 <= heap_bh30_w149_4 & heap_bh30_w149_3 & heap_bh30_w149_5;
   CompressorIn_bh30_422_696 <= heap_bh30_w150_0 & heap_bh30_w150_3;
      Compressor_bh30_422: Compressor_23_3
      port map ( R => CompressorOut_bh30_422_422,
                 X0 => CompressorIn_bh30_422_695,
                 X1 => CompressorIn_bh30_422_696);
   heap_bh30_w149_6 <= CompressorOut_bh30_422_422(0); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w150_4 <= CompressorOut_bh30_422_422(1); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w151_5 <= CompressorOut_bh30_422_422(2); -- cycle= 0 cp= 4.50988e-09

   CompressorIn_bh30_423_697 <= heap_bh30_w161_1 & heap_bh30_w161_0 & heap_bh30_w161_2;
   CompressorIn_bh30_423_698 <= heap_bh30_w162_1 & heap_bh30_w162_0;
      Compressor_bh30_423: Compressor_23_3
      port map ( R => CompressorOut_bh30_423_423,
                 X0 => CompressorIn_bh30_423_697,
                 X1 => CompressorIn_bh30_423_698);
   heap_bh30_w161_3 <= CompressorOut_bh30_423_423(0); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w162_2 <= CompressorOut_bh30_423_423(1); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w163_1 <= CompressorOut_bh30_423_423(2); -- cycle= 0 cp= 4.50988e-09

   CompressorIn_bh30_424_699 <= heap_bh30_w18_11 & heap_bh30_w18_10 & heap_bh30_w18_12;
   CompressorIn_bh30_424_700(0) <= heap_bh30_w19_11;
      Compressor_bh30_424: Compressor_13_3
      port map ( R => CompressorOut_bh30_424_424,
                 X0 => CompressorIn_bh30_424_699,
                 X1 => CompressorIn_bh30_424_700);
   heap_bh30_w18_13 <= CompressorOut_bh30_424_424(0); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w19_12 <= CompressorOut_bh30_424_424(1); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w20_12 <= CompressorOut_bh30_424_424(2); -- cycle= 0 cp= 4.50988e-09

   CompressorIn_bh30_425_701 <= heap_bh30_w26_10 & heap_bh30_w26_13 & heap_bh30_w26_14;
   CompressorIn_bh30_425_702(0) <= heap_bh30_w27_14;
      Compressor_bh30_425: Compressor_13_3
      port map ( R => CompressorOut_bh30_425_425,
                 X0 => CompressorIn_bh30_425_701,
                 X1 => CompressorIn_bh30_425_702);
   heap_bh30_w26_15 <= CompressorOut_bh30_425_425(0); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w27_15 <= CompressorOut_bh30_425_425(1); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w28_16 <= CompressorOut_bh30_425_425(2); -- cycle= 0 cp= 4.50988e-09

   CompressorIn_bh30_426_703 <= heap_bh30_w29_10 & heap_bh30_w29_13 & heap_bh30_w29_14;
   CompressorIn_bh30_426_704(0) <= heap_bh30_w30_14;
      Compressor_bh30_426: Compressor_13_3
      port map ( R => CompressorOut_bh30_426_426,
                 X0 => CompressorIn_bh30_426_703,
                 X1 => CompressorIn_bh30_426_704);
   heap_bh30_w29_15 <= CompressorOut_bh30_426_426(0); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w30_15 <= CompressorOut_bh30_426_426(1); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w31_16 <= CompressorOut_bh30_426_426(2); -- cycle= 0 cp= 4.50988e-09

   CompressorIn_bh30_427_705 <= heap_bh30_w32_10 & heap_bh30_w32_13 & heap_bh30_w32_14;
   CompressorIn_bh30_427_706(0) <= heap_bh30_w33_15;
      Compressor_bh30_427: Compressor_13_3
      port map ( R => CompressorOut_bh30_427_427,
                 X0 => CompressorIn_bh30_427_705,
                 X1 => CompressorIn_bh30_427_706);
   heap_bh30_w32_15 <= CompressorOut_bh30_427_427(0); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w33_16 <= CompressorOut_bh30_427_427(1); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w34_17 <= CompressorOut_bh30_427_427(2); -- cycle= 0 cp= 4.50988e-09

   CompressorIn_bh30_428_707 <= heap_bh30_w37_16 & heap_bh30_w37_15 & heap_bh30_w37_17;
   CompressorIn_bh30_428_708(0) <= heap_bh30_w38_15;
      Compressor_bh30_428: Compressor_13_3
      port map ( R => CompressorOut_bh30_428_428,
                 X0 => CompressorIn_bh30_428_707,
                 X1 => CompressorIn_bh30_428_708);
   heap_bh30_w37_18 <= CompressorOut_bh30_428_428(0); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w38_16 <= CompressorOut_bh30_428_428(1); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w39_18 <= CompressorOut_bh30_428_428(2); -- cycle= 0 cp= 4.50988e-09

   CompressorIn_bh30_429_709 <= heap_bh30_w40_16 & heap_bh30_w40_15 & heap_bh30_w40_17;
   CompressorIn_bh30_429_710(0) <= heap_bh30_w41_15;
      Compressor_bh30_429: Compressor_13_3
      port map ( R => CompressorOut_bh30_429_429,
                 X0 => CompressorIn_bh30_429_709,
                 X1 => CompressorIn_bh30_429_710);
   heap_bh30_w40_18 <= CompressorOut_bh30_429_429(0); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w41_16 <= CompressorOut_bh30_429_429(1); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w42_18 <= CompressorOut_bh30_429_429(2); -- cycle= 0 cp= 4.50988e-09

   CompressorIn_bh30_430_711 <= heap_bh30_w43_16 & heap_bh30_w43_15 & heap_bh30_w43_17;
   CompressorIn_bh30_430_712(0) <= heap_bh30_w44_15;
      Compressor_bh30_430: Compressor_13_3
      port map ( R => CompressorOut_bh30_430_430,
                 X0 => CompressorIn_bh30_430_711,
                 X1 => CompressorIn_bh30_430_712);
   heap_bh30_w43_18 <= CompressorOut_bh30_430_430(0); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w44_16 <= CompressorOut_bh30_430_430(1); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w45_18 <= CompressorOut_bh30_430_430(2); -- cycle= 0 cp= 4.50988e-09

   CompressorIn_bh30_431_713 <= heap_bh30_w51_18 & heap_bh30_w51_17 & heap_bh30_w51_19;
   CompressorIn_bh30_431_714(0) <= heap_bh30_w52_20;
      Compressor_bh30_431: Compressor_13_3
      port map ( R => CompressorOut_bh30_431_431,
                 X0 => CompressorIn_bh30_431_713,
                 X1 => CompressorIn_bh30_431_714);
   heap_bh30_w51_20 <= CompressorOut_bh30_431_431(0); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w52_21 <= CompressorOut_bh30_431_431(1); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w53_20 <= CompressorOut_bh30_431_431(2); -- cycle= 0 cp= 4.50988e-09

   CompressorIn_bh30_432_715 <= heap_bh30_w54_18 & heap_bh30_w54_17 & heap_bh30_w54_19;
   CompressorIn_bh30_432_716(0) <= heap_bh30_w55_20;
      Compressor_bh30_432: Compressor_13_3
      port map ( R => CompressorOut_bh30_432_432,
                 X0 => CompressorIn_bh30_432_715,
                 X1 => CompressorIn_bh30_432_716);
   heap_bh30_w54_20 <= CompressorOut_bh30_432_432(0); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w55_21 <= CompressorOut_bh30_432_432(1); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w56_20 <= CompressorOut_bh30_432_432(2); -- cycle= 0 cp= 4.50988e-09

   CompressorIn_bh30_433_717 <= heap_bh30_w57_18 & heap_bh30_w57_17 & heap_bh30_w57_19;
   CompressorIn_bh30_433_718(0) <= heap_bh30_w58_20;
      Compressor_bh30_433: Compressor_13_3
      port map ( R => CompressorOut_bh30_433_433,
                 X0 => CompressorIn_bh30_433_717,
                 X1 => CompressorIn_bh30_433_718);
   heap_bh30_w57_20 <= CompressorOut_bh30_433_433(0); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w58_21 <= CompressorOut_bh30_433_433(1); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w59_20 <= CompressorOut_bh30_433_433(2); -- cycle= 0 cp= 4.50988e-09

   CompressorIn_bh30_434_719 <= heap_bh30_w60_18 & heap_bh30_w60_17 & heap_bh30_w60_19;
   CompressorIn_bh30_434_720(0) <= heap_bh30_w61_20;
      Compressor_bh30_434: Compressor_13_3
      port map ( R => CompressorOut_bh30_434_434,
                 X0 => CompressorIn_bh30_434_719,
                 X1 => CompressorIn_bh30_434_720);
   heap_bh30_w60_20 <= CompressorOut_bh30_434_434(0); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w61_21 <= CompressorOut_bh30_434_434(1); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w62_20 <= CompressorOut_bh30_434_434(2); -- cycle= 0 cp= 4.50988e-09

   CompressorIn_bh30_435_721 <= heap_bh30_w63_18 & heap_bh30_w63_17 & heap_bh30_w63_19;
   CompressorIn_bh30_435_722(0) <= heap_bh30_w64_20;
      Compressor_bh30_435: Compressor_13_3
      port map ( R => CompressorOut_bh30_435_435,
                 X0 => CompressorIn_bh30_435_721,
                 X1 => CompressorIn_bh30_435_722);
   heap_bh30_w63_20 <= CompressorOut_bh30_435_435(0); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w64_21 <= CompressorOut_bh30_435_435(1); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w65_20 <= CompressorOut_bh30_435_435(2); -- cycle= 0 cp= 4.50988e-09

   CompressorIn_bh30_436_723 <= heap_bh30_w66_18 & heap_bh30_w66_17 & heap_bh30_w66_19;
   CompressorIn_bh30_436_724(0) <= heap_bh30_w67_21;
      Compressor_bh30_436: Compressor_13_3
      port map ( R => CompressorOut_bh30_436_436,
                 X0 => CompressorIn_bh30_436_723,
                 X1 => CompressorIn_bh30_436_724);
   heap_bh30_w66_20 <= CompressorOut_bh30_436_436(0); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w67_22 <= CompressorOut_bh30_436_436(1); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w68_21 <= CompressorOut_bh30_436_436(2); -- cycle= 0 cp= 4.50988e-09

   CompressorIn_bh30_437_725 <= heap_bh30_w71_21 & heap_bh30_w71_20 & heap_bh30_w71_22;
   CompressorIn_bh30_437_726(0) <= heap_bh30_w72_24;
      Compressor_bh30_437: Compressor_13_3
      port map ( R => CompressorOut_bh30_437_437,
                 X0 => CompressorIn_bh30_437_725,
                 X1 => CompressorIn_bh30_437_726);
   heap_bh30_w71_23 <= CompressorOut_bh30_437_437(0); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w72_25 <= CompressorOut_bh30_437_437(1); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w73_24 <= CompressorOut_bh30_437_437(2); -- cycle= 0 cp= 4.50988e-09

   CompressorIn_bh30_438_727 <= heap_bh30_w110_11 & heap_bh30_w110_10 & heap_bh30_w110_12;
   CompressorIn_bh30_438_728(0) <= heap_bh30_w111_13;
      Compressor_bh30_438: Compressor_13_3
      port map ( R => CompressorOut_bh30_438_438,
                 X0 => CompressorIn_bh30_438_727,
                 X1 => CompressorIn_bh30_438_728);
   heap_bh30_w110_13 <= CompressorOut_bh30_438_438(0); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w111_14 <= CompressorOut_bh30_438_438(1); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w112_11 <= CompressorOut_bh30_438_438(2); -- cycle= 0 cp= 4.50988e-09

   CompressorIn_bh30_439_729 <= heap_bh30_w68_17 & heap_bh30_w68_20 & heap_bh30_w68_21;
   CompressorIn_bh30_439_730 <= heap_bh30_w69_23 & heap_bh30_w69_22;
      Compressor_bh30_439: Compressor_23_3
      port map ( R => CompressorOut_bh30_439_439,
                 X0 => CompressorIn_bh30_439_729,
                 X1 => CompressorIn_bh30_439_730);
   heap_bh30_w68_22 <= CompressorOut_bh30_439_439(0); -- cycle= 0 cp= 5.0406e-09
   heap_bh30_w69_24 <= CompressorOut_bh30_439_439(1); -- cycle= 0 cp= 5.0406e-09
   heap_bh30_w70_23 <= CompressorOut_bh30_439_439(2); -- cycle= 0 cp= 5.0406e-09

   CompressorIn_bh30_440_731 <= heap_bh30_w73_20 & heap_bh30_w73_23 & heap_bh30_w73_24;
   CompressorIn_bh30_440_732 <= heap_bh30_w74_24 & heap_bh30_w74_23;
      Compressor_bh30_440: Compressor_23_3
      port map ( R => CompressorOut_bh30_440_440,
                 X0 => CompressorIn_bh30_440_731,
                 X1 => CompressorIn_bh30_440_732);
   heap_bh30_w73_25 <= CompressorOut_bh30_440_440(0); -- cycle= 0 cp= 5.0406e-09
   heap_bh30_w74_25 <= CompressorOut_bh30_440_440(1); -- cycle= 0 cp= 5.0406e-09
   heap_bh30_w75_26 <= CompressorOut_bh30_440_440(2); -- cycle= 0 cp= 5.0406e-09

   CompressorIn_bh30_441_733 <= heap_bh30_w95_12 & heap_bh30_w95_15 & heap_bh30_w95_16;
   CompressorIn_bh30_441_734 <= heap_bh30_w96_15 & heap_bh30_w96_14;
      Compressor_bh30_441: Compressor_23_3
      port map ( R => CompressorOut_bh30_441_441,
                 X0 => CompressorIn_bh30_441_733,
                 X1 => CompressorIn_bh30_441_734);
   heap_bh30_w95_17 <= CompressorOut_bh30_441_441(0); -- cycle= 0 cp= 5.0406e-09
   heap_bh30_w96_16 <= CompressorOut_bh30_441_441(1); -- cycle= 0 cp= 5.0406e-09
   heap_bh30_w97_16 <= CompressorOut_bh30_441_441(2); -- cycle= 0 cp= 5.0406e-09

   CompressorIn_bh30_442_735 <= heap_bh30_w99_11 & heap_bh30_w99_14 & heap_bh30_w99_15;
   CompressorIn_bh30_442_736 <= heap_bh30_w100_15 & heap_bh30_w100_14;
      Compressor_bh30_442: Compressor_23_3
      port map ( R => CompressorOut_bh30_442_442,
                 X0 => CompressorIn_bh30_442_735,
                 X1 => CompressorIn_bh30_442_736);
   heap_bh30_w99_16 <= CompressorOut_bh30_442_442(0); -- cycle= 0 cp= 5.0406e-09
   heap_bh30_w100_16 <= CompressorOut_bh30_442_442(1); -- cycle= 0 cp= 5.0406e-09
   heap_bh30_w101_15 <= CompressorOut_bh30_442_442(2); -- cycle= 0 cp= 5.0406e-09

   CompressorIn_bh30_443_737 <= heap_bh30_w115_10 & heap_bh30_w115_9 & heap_bh30_w115_11;
   CompressorIn_bh30_443_738 <= heap_bh30_w116_6 & heap_bh30_w116_9;
      Compressor_bh30_443: Compressor_23_3
      port map ( R => CompressorOut_bh30_443_443,
                 X0 => CompressorIn_bh30_443_737,
                 X1 => CompressorIn_bh30_443_738);
   heap_bh30_w115_12 <= CompressorOut_bh30_443_443(0); -- cycle= 0 cp= 5.0406e-09
   heap_bh30_w116_10 <= CompressorOut_bh30_443_443(1); -- cycle= 0 cp= 5.0406e-09
   heap_bh30_w117_11 <= CompressorOut_bh30_443_443(2); -- cycle= 0 cp= 5.0406e-09

   CompressorIn_bh30_444_739 <= heap_bh30_w151_4 & heap_bh30_w151_3 & heap_bh30_w151_5;
   CompressorIn_bh30_444_740 <= heap_bh30_w152_0 & heap_bh30_w152_3;
      Compressor_bh30_444: Compressor_23_3
      port map ( R => CompressorOut_bh30_444_444,
                 X0 => CompressorIn_bh30_444_739,
                 X1 => CompressorIn_bh30_444_740);
   heap_bh30_w151_6 <= CompressorOut_bh30_444_444(0); -- cycle= 0 cp= 5.0406e-09
   heap_bh30_w152_4 <= CompressorOut_bh30_444_444(1); -- cycle= 0 cp= 5.0406e-09
   heap_bh30_w153_5 <= CompressorOut_bh30_444_444(2); -- cycle= 0 cp= 5.0406e-09

   CompressorIn_bh30_445_741 <= heap_bh30_w48_17 & heap_bh30_w48_16 & heap_bh30_w48_18;
   CompressorIn_bh30_445_742(0) <= heap_bh30_w49_17;
      Compressor_bh30_445: Compressor_13_3
      port map ( R => CompressorOut_bh30_445_445,
                 X0 => CompressorIn_bh30_445_741,
                 X1 => CompressorIn_bh30_445_742);
   heap_bh30_w48_19 <= CompressorOut_bh30_445_445(0); -- cycle= 0 cp= 5.0406e-09
   heap_bh30_w49_18 <= CompressorOut_bh30_445_445(1); -- cycle= 0 cp= 5.0406e-09
   heap_bh30_w50_19 <= CompressorOut_bh30_445_445(2); -- cycle= 0 cp= 5.0406e-09

   CompressorIn_bh30_446_743 <= heap_bh30_w53_16 & heap_bh30_w53_19 & heap_bh30_w53_20;
   CompressorIn_bh30_446_744(0) <= heap_bh30_w54_20;
      Compressor_bh30_446: Compressor_13_3
      port map ( R => CompressorOut_bh30_446_446,
                 X0 => CompressorIn_bh30_446_743,
                 X1 => CompressorIn_bh30_446_744);
   heap_bh30_w53_21 <= CompressorOut_bh30_446_446(0); -- cycle= 0 cp= 5.0406e-09
   heap_bh30_w54_21 <= CompressorOut_bh30_446_446(1); -- cycle= 0 cp= 5.0406e-09
   heap_bh30_w55_22 <= CompressorOut_bh30_446_446(2); -- cycle= 0 cp= 5.0406e-09

   CompressorIn_bh30_447_745 <= heap_bh30_w56_16 & heap_bh30_w56_19 & heap_bh30_w56_20;
   CompressorIn_bh30_447_746(0) <= heap_bh30_w57_20;
      Compressor_bh30_447: Compressor_13_3
      port map ( R => CompressorOut_bh30_447_447,
                 X0 => CompressorIn_bh30_447_745,
                 X1 => CompressorIn_bh30_447_746);
   heap_bh30_w56_21 <= CompressorOut_bh30_447_447(0); -- cycle= 0 cp= 5.0406e-09
   heap_bh30_w57_21 <= CompressorOut_bh30_447_447(1); -- cycle= 0 cp= 5.0406e-09
   heap_bh30_w58_22 <= CompressorOut_bh30_447_447(2); -- cycle= 0 cp= 5.0406e-09

   CompressorIn_bh30_448_747 <= heap_bh30_w59_16 & heap_bh30_w59_19 & heap_bh30_w59_20;
   CompressorIn_bh30_448_748(0) <= heap_bh30_w60_20;
      Compressor_bh30_448: Compressor_13_3
      port map ( R => CompressorOut_bh30_448_448,
                 X0 => CompressorIn_bh30_448_747,
                 X1 => CompressorIn_bh30_448_748);
   heap_bh30_w59_21 <= CompressorOut_bh30_448_448(0); -- cycle= 0 cp= 5.0406e-09
   heap_bh30_w60_21 <= CompressorOut_bh30_448_448(1); -- cycle= 0 cp= 5.0406e-09
   heap_bh30_w61_22 <= CompressorOut_bh30_448_448(2); -- cycle= 0 cp= 5.0406e-09

   CompressorIn_bh30_449_749 <= heap_bh30_w62_16 & heap_bh30_w62_19 & heap_bh30_w62_20;
   CompressorIn_bh30_449_750(0) <= heap_bh30_w63_20;
      Compressor_bh30_449: Compressor_13_3
      port map ( R => CompressorOut_bh30_449_449,
                 X0 => CompressorIn_bh30_449_749,
                 X1 => CompressorIn_bh30_449_750);
   heap_bh30_w62_21 <= CompressorOut_bh30_449_449(0); -- cycle= 0 cp= 5.0406e-09
   heap_bh30_w63_21 <= CompressorOut_bh30_449_449(1); -- cycle= 0 cp= 5.0406e-09
   heap_bh30_w64_22 <= CompressorOut_bh30_449_449(2); -- cycle= 0 cp= 5.0406e-09

   CompressorIn_bh30_450_751 <= heap_bh30_w65_16 & heap_bh30_w65_19 & heap_bh30_w65_20;
   CompressorIn_bh30_450_752(0) <= heap_bh30_w66_20;
      Compressor_bh30_450: Compressor_13_3
      port map ( R => CompressorOut_bh30_450_450,
                 X0 => CompressorIn_bh30_450_751,
                 X1 => CompressorIn_bh30_450_752);
   heap_bh30_w65_21 <= CompressorOut_bh30_450_450(0); -- cycle= 0 cp= 5.0406e-09
   heap_bh30_w66_21 <= CompressorOut_bh30_450_450(1); -- cycle= 0 cp= 5.0406e-09
   heap_bh30_w67_23 <= CompressorOut_bh30_450_450(2); -- cycle= 0 cp= 5.0406e-09

   CompressorIn_bh30_451_753 <= heap_bh30_w77_24 & heap_bh30_w77_23 & heap_bh30_w77_25;
   CompressorIn_bh30_451_754(0) <= heap_bh30_w78_25;
      Compressor_bh30_451: Compressor_13_3
      port map ( R => CompressorOut_bh30_451_451,
                 X0 => CompressorIn_bh30_451_753,
                 X1 => CompressorIn_bh30_451_754);
   heap_bh30_w77_26 <= CompressorOut_bh30_451_451(0); -- cycle= 0 cp= 5.0406e-09
   heap_bh30_w78_26 <= CompressorOut_bh30_451_451(1); -- cycle= 0 cp= 5.0406e-09
   heap_bh30_w79_26 <= CompressorOut_bh30_451_451(2); -- cycle= 0 cp= 5.0406e-09

   CompressorIn_bh30_452_755 <= heap_bh30_w80_24 & heap_bh30_w80_23 & heap_bh30_w80_25;
   CompressorIn_bh30_452_756(0) <= heap_bh30_w81_25;
      Compressor_bh30_452: Compressor_13_3
      port map ( R => CompressorOut_bh30_452_452,
                 X0 => CompressorIn_bh30_452_755,
                 X1 => CompressorIn_bh30_452_756);
   heap_bh30_w80_26 <= CompressorOut_bh30_452_452(0); -- cycle= 0 cp= 5.0406e-09
   heap_bh30_w81_26 <= CompressorOut_bh30_452_452(1); -- cycle= 0 cp= 5.0406e-09
   heap_bh30_w82_26 <= CompressorOut_bh30_452_452(2); -- cycle= 0 cp= 5.0406e-09

   CompressorIn_bh30_453_757 <= heap_bh30_w83_24 & heap_bh30_w83_23 & heap_bh30_w83_25;
   CompressorIn_bh30_453_758(0) <= heap_bh30_w84_25;
      Compressor_bh30_453: Compressor_13_3
      port map ( R => CompressorOut_bh30_453_453,
                 X0 => CompressorIn_bh30_453_757,
                 X1 => CompressorIn_bh30_453_758);
   heap_bh30_w83_26 <= CompressorOut_bh30_453_453(0); -- cycle= 0 cp= 5.0406e-09
   heap_bh30_w84_26 <= CompressorOut_bh30_453_453(1); -- cycle= 0 cp= 5.0406e-09
   heap_bh30_w85_26 <= CompressorOut_bh30_453_453(2); -- cycle= 0 cp= 5.0406e-09

   CompressorIn_bh30_454_759 <= heap_bh30_w86_24 & heap_bh30_w86_23 & heap_bh30_w86_25;
   CompressorIn_bh30_454_760(0) <= heap_bh30_w87_25;
      Compressor_bh30_454: Compressor_13_3
      port map ( R => CompressorOut_bh30_454_454,
                 X0 => CompressorIn_bh30_454_759,
                 X1 => CompressorIn_bh30_454_760);
   heap_bh30_w86_26 <= CompressorOut_bh30_454_454(0); -- cycle= 0 cp= 5.0406e-09
   heap_bh30_w87_26 <= CompressorOut_bh30_454_454(1); -- cycle= 0 cp= 5.0406e-09
   heap_bh30_w88_26 <= CompressorOut_bh30_454_454(2); -- cycle= 0 cp= 5.0406e-09

   CompressorIn_bh30_455_761 <= heap_bh30_w89_24 & heap_bh30_w89_23 & heap_bh30_w89_25;
   CompressorIn_bh30_455_762(0) <= heap_bh30_w90_24;
      Compressor_bh30_455: Compressor_13_3
      port map ( R => CompressorOut_bh30_455_455,
                 X0 => CompressorIn_bh30_455_761,
                 X1 => CompressorIn_bh30_455_762);
   heap_bh30_w89_26 <= CompressorOut_bh30_455_455(0); -- cycle= 0 cp= 5.0406e-09
   heap_bh30_w90_25 <= CompressorOut_bh30_455_455(1); -- cycle= 0 cp= 5.0406e-09
   heap_bh30_w91_24 <= CompressorOut_bh30_455_455(2); -- cycle= 0 cp= 5.0406e-09

   CompressorIn_bh30_456_763 <= heap_bh30_w92_20 & heap_bh30_w92_19 & heap_bh30_w92_21;
   CompressorIn_bh30_456_764(0) <= heap_bh30_w93_19;
      Compressor_bh30_456: Compressor_13_3
      port map ( R => CompressorOut_bh30_456_456,
                 X0 => CompressorIn_bh30_456_763,
                 X1 => CompressorIn_bh30_456_764);
   heap_bh30_w92_22 <= CompressorOut_bh30_456_456(0); -- cycle= 0 cp= 5.0406e-09
   heap_bh30_w93_20 <= CompressorOut_bh30_456_456(1); -- cycle= 0 cp= 5.0406e-09
   heap_bh30_w94_19 <= CompressorOut_bh30_456_456(2); -- cycle= 0 cp= 5.0406e-09

   CompressorIn_bh30_457_765 <= heap_bh30_w112_9 & heap_bh30_w112_10 & heap_bh30_w112_11;
   CompressorIn_bh30_457_766(0) <= heap_bh30_w113_12;
      Compressor_bh30_457: Compressor_13_3
      port map ( R => CompressorOut_bh30_457_457,
                 X0 => CompressorIn_bh30_457_765,
                 X1 => CompressorIn_bh30_457_766);
   heap_bh30_w112_12 <= CompressorOut_bh30_457_457(0); -- cycle= 0 cp= 5.0406e-09
   heap_bh30_w113_13 <= CompressorOut_bh30_457_457(1); -- cycle= 0 cp= 5.0406e-09
   heap_bh30_w114_11 <= CompressorOut_bh30_457_457(2); -- cycle= 0 cp= 5.0406e-09

   CompressorIn_bh30_458_767 <= heap_bh30_w101_11 & heap_bh30_w101_14 & heap_bh30_w101_15;
   CompressorIn_bh30_458_768 <= heap_bh30_w102_15 & heap_bh30_w102_14;
      Compressor_bh30_458: Compressor_23_3
      port map ( R => CompressorOut_bh30_458_458,
                 X0 => CompressorIn_bh30_458_767,
                 X1 => CompressorIn_bh30_458_768);
   heap_bh30_w101_16 <= CompressorOut_bh30_458_458(0); -- cycle= 0 cp= 5.57132e-09
   heap_bh30_w102_16 <= CompressorOut_bh30_458_458(1); -- cycle= 0 cp= 5.57132e-09
   heap_bh30_w103_15 <= CompressorOut_bh30_458_458(2); -- cycle= 0 cp= 5.57132e-09

   CompressorIn_bh30_459_769 <= heap_bh30_w117_10 & heap_bh30_w117_9 & heap_bh30_w117_11;
   CompressorIn_bh30_459_770 <= heap_bh30_w118_6 & heap_bh30_w118_9;
      Compressor_bh30_459: Compressor_23_3
      port map ( R => CompressorOut_bh30_459_459,
                 X0 => CompressorIn_bh30_459_769,
                 X1 => CompressorIn_bh30_459_770);
   heap_bh30_w117_12 <= CompressorOut_bh30_459_459(0); -- cycle= 0 cp= 5.57132e-09
   heap_bh30_w118_10 <= CompressorOut_bh30_459_459(1); -- cycle= 0 cp= 5.57132e-09
   heap_bh30_w119_11 <= CompressorOut_bh30_459_459(2); -- cycle= 0 cp= 5.57132e-09

   CompressorIn_bh30_460_771 <= heap_bh30_w153_4 & heap_bh30_w153_3 & heap_bh30_w153_5;
   CompressorIn_bh30_460_772 <= heap_bh30_w154_0 & heap_bh30_w154_3;
      Compressor_bh30_460: Compressor_23_3
      port map ( R => CompressorOut_bh30_460_460,
                 X0 => CompressorIn_bh30_460_771,
                 X1 => CompressorIn_bh30_460_772);
   heap_bh30_w153_6 <= CompressorOut_bh30_460_460(0); -- cycle= 0 cp= 5.57132e-09
   heap_bh30_w154_4 <= CompressorOut_bh30_460_460(1); -- cycle= 0 cp= 5.57132e-09
   heap_bh30_w155_5 <= CompressorOut_bh30_460_460(2); -- cycle= 0 cp= 5.57132e-09

   CompressorIn_bh30_461_773 <= heap_bh30_w70_19 & heap_bh30_w70_22 & heap_bh30_w70_23;
   CompressorIn_bh30_461_774(0) <= heap_bh30_w71_23;
      Compressor_bh30_461: Compressor_13_3
      port map ( R => CompressorOut_bh30_461_461,
                 X0 => CompressorIn_bh30_461_773,
                 X1 => CompressorIn_bh30_461_774);
   heap_bh30_w70_24 <= CompressorOut_bh30_461_461(0); -- cycle= 0 cp= 5.57132e-09
   heap_bh30_w71_24 <= CompressorOut_bh30_461_461(1); -- cycle= 0 cp= 5.57132e-09
   heap_bh30_w72_26 <= CompressorOut_bh30_461_461(2); -- cycle= 0 cp= 5.57132e-09

   CompressorIn_bh30_462_775 <= heap_bh30_w103_11 & heap_bh30_w103_14 & heap_bh30_w103_15;
   CompressorIn_bh30_462_776 <= heap_bh30_w104_15 & heap_bh30_w104_14;
      Compressor_bh30_462: Compressor_23_3
      port map ( R => CompressorOut_bh30_462_462,
                 X0 => CompressorIn_bh30_462_775,
                 X1 => CompressorIn_bh30_462_776);
   heap_bh30_w103_16 <= CompressorOut_bh30_462_462(0); -- cycle= 0 cp= 6.10204e-09
   heap_bh30_w104_16 <= CompressorOut_bh30_462_462(1); -- cycle= 0 cp= 6.10204e-09
   heap_bh30_w105_15 <= CompressorOut_bh30_462_462(2); -- cycle= 0 cp= 6.10204e-09

   CompressorIn_bh30_463_777 <= heap_bh30_w119_10 & heap_bh30_w119_9 & heap_bh30_w119_11;
   CompressorIn_bh30_463_778 <= heap_bh30_w120_6 & heap_bh30_w120_9;
      Compressor_bh30_463: Compressor_23_3
      port map ( R => CompressorOut_bh30_463_463,
                 X0 => CompressorIn_bh30_463_777,
                 X1 => CompressorIn_bh30_463_778);
   heap_bh30_w119_12 <= CompressorOut_bh30_463_463(0); -- cycle= 0 cp= 6.10204e-09
   heap_bh30_w120_10 <= CompressorOut_bh30_463_463(1); -- cycle= 0 cp= 6.10204e-09
   heap_bh30_w121_11 <= CompressorOut_bh30_463_463(2); -- cycle= 0 cp= 6.10204e-09

   CompressorIn_bh30_464_779 <= heap_bh30_w155_4 & heap_bh30_w155_3 & heap_bh30_w155_5;
   CompressorIn_bh30_464_780(0) <= heap_bh30_w156_2;
      Compressor_bh30_464: Compressor_13_3
      port map ( R => CompressorOut_bh30_464_464,
                 X0 => CompressorIn_bh30_464_779,
                 X1 => CompressorIn_bh30_464_780);
   heap_bh30_w155_6 <= CompressorOut_bh30_464_464(0); -- cycle= 0 cp= 6.10204e-09
   heap_bh30_w156_3 <= CompressorOut_bh30_464_464(1); -- cycle= 0 cp= 6.10204e-09
   heap_bh30_w157_4 <= CompressorOut_bh30_464_464(2); -- cycle= 0 cp= 6.10204e-09

   CompressorIn_bh30_465_781 <= heap_bh30_w105_11 & heap_bh30_w105_14 & heap_bh30_w105_15;
   CompressorIn_bh30_465_782 <= heap_bh30_w106_15 & heap_bh30_w106_14;
      Compressor_bh30_465: Compressor_23_3
      port map ( R => CompressorOut_bh30_465_465,
                 X0 => CompressorIn_bh30_465_781,
                 X1 => CompressorIn_bh30_465_782);
   heap_bh30_w105_16 <= CompressorOut_bh30_465_465(0); -- cycle= 0 cp= 6.63276e-09
   heap_bh30_w106_16 <= CompressorOut_bh30_465_465(1); -- cycle= 0 cp= 6.63276e-09
   heap_bh30_w107_15 <= CompressorOut_bh30_465_465(2); -- cycle= 0 cp= 6.63276e-09

   CompressorIn_bh30_466_783 <= heap_bh30_w121_10 & heap_bh30_w121_9 & heap_bh30_w121_11;
   CompressorIn_bh30_466_784 <= heap_bh30_w122_6 & heap_bh30_w122_9;
      Compressor_bh30_466: Compressor_23_3
      port map ( R => CompressorOut_bh30_466_466,
                 X0 => CompressorIn_bh30_466_783,
                 X1 => CompressorIn_bh30_466_784);
   heap_bh30_w121_12 <= CompressorOut_bh30_466_466(0); -- cycle= 0 cp= 6.63276e-09
   heap_bh30_w122_10 <= CompressorOut_bh30_466_466(1); -- cycle= 0 cp= 6.63276e-09
   heap_bh30_w123_11 <= CompressorOut_bh30_466_466(2); -- cycle= 0 cp= 6.63276e-09

   CompressorIn_bh30_467_785 <= heap_bh30_w107_11 & heap_bh30_w107_14 & heap_bh30_w107_15;
   CompressorIn_bh30_467_786 <= heap_bh30_w108_14 & heap_bh30_w108_13;
      Compressor_bh30_467: Compressor_23_3
      port map ( R => CompressorOut_bh30_467_467,
                 X0 => CompressorIn_bh30_467_785,
                 X1 => CompressorIn_bh30_467_786);
   heap_bh30_w107_16 <= CompressorOut_bh30_467_467(0); -- cycle= 0 cp= 7.16348e-09
   heap_bh30_w108_15 <= CompressorOut_bh30_467_467(1); -- cycle= 0 cp= 7.16348e-09
   heap_bh30_w109_14 <= CompressorOut_bh30_467_467(2); -- cycle= 0 cp= 7.16348e-09

   CompressorIn_bh30_468_787 <= heap_bh30_w123_10 & heap_bh30_w123_9 & heap_bh30_w123_11;
   CompressorIn_bh30_468_788 <= heap_bh30_w124_6 & heap_bh30_w124_9;
      Compressor_bh30_468: Compressor_23_3
      port map ( R => CompressorOut_bh30_468_468,
                 X0 => CompressorIn_bh30_468_787,
                 X1 => CompressorIn_bh30_468_788);
   heap_bh30_w123_12 <= CompressorOut_bh30_468_468(0); -- cycle= 0 cp= 7.16348e-09
   heap_bh30_w124_10 <= CompressorOut_bh30_468_468(1); -- cycle= 0 cp= 7.16348e-09
   heap_bh30_w125_11 <= CompressorOut_bh30_468_468(2); -- cycle= 0 cp= 7.16348e-09

   CompressorIn_bh30_469_789 <= heap_bh30_w125_10 & heap_bh30_w125_9 & heap_bh30_w125_11;
   CompressorIn_bh30_469_790 <= heap_bh30_w126_6 & heap_bh30_w126_9;
      Compressor_bh30_469: Compressor_23_3
      port map ( R => CompressorOut_bh30_469_469,
                 X0 => CompressorIn_bh30_469_789,
                 X1 => CompressorIn_bh30_469_790);
   heap_bh30_w125_12 <= CompressorOut_bh30_469_469(0); -- cycle= 0 cp= 7.6942e-09
   heap_bh30_w126_10 <= CompressorOut_bh30_469_469(1); -- cycle= 0 cp= 7.6942e-09
   heap_bh30_w127_11 <= CompressorOut_bh30_469_469(2); -- cycle= 0 cp= 7.6942e-09

   CompressorIn_bh30_470_791 <= heap_bh30_w109_10 & heap_bh30_w109_13 & heap_bh30_w109_14;
   CompressorIn_bh30_470_792(0) <= heap_bh30_w110_13;
      Compressor_bh30_470: Compressor_13_3
      port map ( R => CompressorOut_bh30_470_470,
                 X0 => CompressorIn_bh30_470_791,
                 X1 => CompressorIn_bh30_470_792);
   heap_bh30_w109_15 <= CompressorOut_bh30_470_470(0); -- cycle= 0 cp= 7.6942e-09
   heap_bh30_w110_14 <= CompressorOut_bh30_470_470(1); -- cycle= 0 cp= 7.6942e-09
   heap_bh30_w111_15 <= CompressorOut_bh30_470_470(2); -- cycle= 0 cp= 7.6942e-09

   CompressorIn_bh30_471_793 <= heap_bh30_w127_10 & heap_bh30_w127_9 & heap_bh30_w127_11;
   CompressorIn_bh30_471_794 <= heap_bh30_w128_6 & heap_bh30_w128_9;
      Compressor_bh30_471: Compressor_23_3
      port map ( R => CompressorOut_bh30_471_471,
                 X0 => CompressorIn_bh30_471_793,
                 X1 => CompressorIn_bh30_471_794);
   heap_bh30_w127_12 <= CompressorOut_bh30_471_471(0); -- cycle= 0 cp= 8.22492e-09
   heap_bh30_w128_10 <= CompressorOut_bh30_471_471(1); -- cycle= 0 cp= 8.22492e-09
   heap_bh30_w129_10 <= CompressorOut_bh30_471_471(2); -- cycle= 0 cp= 8.22492e-09

   CompressorIn_bh30_472_795 <= heap_bh30_w129_9 & heap_bh30_w129_8 & heap_bh30_w129_10;
   CompressorIn_bh30_472_796(0) <= heap_bh30_w130_9;
      Compressor_bh30_472: Compressor_13_3
      port map ( R => CompressorOut_bh30_472_472,
                 X0 => CompressorIn_bh30_472_795,
                 X1 => CompressorIn_bh30_472_796);
   heap_bh30_w129_11 <= CompressorOut_bh30_472_472(0); -- cycle= 0 cp= 8.75564e-09
   heap_bh30_w130_10 <= CompressorOut_bh30_472_472(1); -- cycle= 0 cp= 8.75564e-09
   heap_bh30_w131_11 <= CompressorOut_bh30_472_472(2); -- cycle= 0 cp= 8.75564e-09
   finalAdderIn0_bh30 <= "0" & heap_bh30_w179_0 & heap_bh30_w178_0 & heap_bh30_w177_0 & heap_bh30_w176_0 & heap_bh30_w175_0 & heap_bh30_w174_0 & heap_bh30_w173_0 & heap_bh30_w172_0 & heap_bh30_w171_0 & heap_bh30_w170_0 & heap_bh30_w169_0 & heap_bh30_w168_0 & heap_bh30_w167_0 & heap_bh30_w166_0 & heap_bh30_w165_0 & heap_bh30_w164_0 & heap_bh30_w163_0 & heap_bh30_w162_2 & heap_bh30_w161_3 & heap_bh30_w160_2 & heap_bh30_w159_3 & heap_bh30_w158_2 & heap_bh30_w157_3 & heap_bh30_w156_3 & heap_bh30_w155_6 & heap_bh30_w154_4 & heap_bh30_w153_6 & heap_bh30_w152_4 & heap_bh30_w151_6 & heap_bh30_w150_4 & heap_bh30_w149_6 & heap_bh30_w148_4 & heap_bh30_w147_6 & heap_bh30_w146_3 & heap_bh30_w145_8 & heap_bh30_w144_6 & heap_bh30_w143_8 & heap_bh30_w142_6 & heap_bh30_w141_8 & heap_bh30_w140_6 & heap_bh30_w139_8 & heap_bh30_w138_6 & heap_bh30_w137_8 & heap_bh30_w136_6 & heap_bh30_w135_8 & heap_bh30_w134_6 & heap_bh30_w133_9 & heap_bh30_w132_9 & heap_bh30_w131_10 & heap_bh30_w130_10 & heap_bh30_w129_11 & heap_bh30_w128_10 & heap_bh30_w127_12 & heap_bh30_w126_10 & heap_bh30_w125_12 & heap_bh30_w124_10 & heap_bh30_w123_12 & heap_bh30_w122_10 & heap_bh30_w121_12 & heap_bh30_w120_10 & heap_bh30_w119_12 & heap_bh30_w118_10 & heap_bh30_w117_12 & heap_bh30_w116_10 & heap_bh30_w115_12 & heap_bh30_w114_10 & heap_bh30_w113_13 & heap_bh30_w112_12 & heap_bh30_w111_14 & heap_bh30_w110_14 & heap_bh30_w109_15 & heap_bh30_w108_15 & heap_bh30_w107_16 & heap_bh30_w106_16 & heap_bh30_w105_16 & heap_bh30_w104_16 & heap_bh30_w103_16 & heap_bh30_w102_16 & heap_bh30_w101_16 & heap_bh30_w100_16 & heap_bh30_w99_16 & heap_bh30_w98_16 & heap_bh30_w97_15 & heap_bh30_w96_16 & heap_bh30_w95_17 & heap_bh30_w94_18 & heap_bh30_w93_20 & heap_bh30_w92_22 & heap_bh30_w91_23 & heap_bh30_w90_25 & heap_bh30_w89_26 & heap_bh30_w88_25 & heap_bh30_w87_26 & heap_bh30_w86_26 & heap_bh30_w85_25 & heap_bh30_w84_26 & heap_bh30_w83_26 & heap_bh30_w82_25 & heap_bh30_w81_26 & heap_bh30_w80_26 & heap_bh30_w79_25 & heap_bh30_w78_26 & heap_bh30_w77_26 & heap_bh30_w76_25 & heap_bh30_w75_25 & heap_bh30_w74_25 & heap_bh30_w73_25 & heap_bh30_w72_25 & heap_bh30_w71_24 & heap_bh30_w70_24 & heap_bh30_w69_24 & heap_bh30_w68_22 & heap_bh30_w67_22 & heap_bh30_w66_21 & heap_bh30_w65_21 & heap_bh30_w64_21 & heap_bh30_w63_21 & heap_bh30_w62_21 & heap_bh30_w61_21 & heap_bh30_w60_21 & heap_bh30_w59_21 & heap_bh30_w58_21 & heap_bh30_w57_21 & heap_bh30_w56_21 & heap_bh30_w55_21 & heap_bh30_w54_21 & heap_bh30_w53_21 & heap_bh30_w52_21 & heap_bh30_w51_20 & heap_bh30_w50_18 & heap_bh30_w49_18 & heap_bh30_w48_19 & heap_bh30_w47_17 & heap_bh30_w46_17 & heap_bh30_w45_17 & heap_bh30_w44_16 & heap_bh30_w43_18 & heap_bh30_w42_17 & heap_bh30_w41_16 & heap_bh30_w40_18 & heap_bh30_w39_17 & heap_bh30_w38_16 & heap_bh30_w37_18 & heap_bh30_w36_17 & heap_bh30_w35_16 & heap_bh30_w34_16 & heap_bh30_w33_16 & heap_bh30_w32_15 & heap_bh30_w31_15 & heap_bh30_w30_15 & heap_bh30_w29_15 & heap_bh30_w28_15 & heap_bh30_w27_15 & heap_bh30_w26_15 & heap_bh30_w25_15 & heap_bh30_w24_14 & heap_bh30_w23_12 & heap_bh30_w22_12 & heap_bh30_w21_13 & heap_bh30_w20_11 & heap_bh30_w19_12 & heap_bh30_w18_13 & heap_bh30_w17_11 & heap_bh30_w16_12 & heap_bh30_w15_10 & heap_bh30_w14_9 & heap_bh30_w13_9 & heap_bh30_w12_9 & heap_bh30_w11_8 & heap_bh30_w10_10 & heap_bh30_w9_8 & heap_bh30_w8_8 & heap_bh30_w7_4 & heap_bh30_w6_8 & heap_bh30_w5_3 & heap_bh30_w4_6 & heap_bh30_w3_5 & heap_bh30_w2_3 & heap_bh30_w1_0 & heap_bh30_w0_0;
   finalAdderIn1_bh30 <= "0" & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & heap_bh30_w163_1 & '0' & '0' & '0' & '0' & '0' & heap_bh30_w157_4 & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & heap_bh30_w146_4 & heap_bh30_w145_7 & '0' & heap_bh30_w143_7 & '0' & heap_bh30_w141_7 & '0' & heap_bh30_w139_7 & '0' & heap_bh30_w137_7 & '0' & heap_bh30_w135_7 & heap_bh30_w134_7 & '0' & '0' & heap_bh30_w131_11 & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & heap_bh30_w114_11 & '0' & '0' & heap_bh30_w111_15 & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & heap_bh30_w97_16 & '0' & '0' & heap_bh30_w94_19 & '0' & '0' & heap_bh30_w91_24 & '0' & '0' & heap_bh30_w88_26 & '0' & '0' & heap_bh30_w85_26 & '0' & '0' & heap_bh30_w82_26 & '0' & '0' & heap_bh30_w79_26 & '0' & '0' & '0' & heap_bh30_w75_26 & '0' & '0' & heap_bh30_w72_26 & '0' & '0' & '0' & '0' & heap_bh30_w67_23 & '0' & '0' & heap_bh30_w64_22 & '0' & '0' & heap_bh30_w61_22 & '0' & '0' & heap_bh30_w58_22 & '0' & '0' & heap_bh30_w55_22 & '0' & '0' & '0' & '0' & heap_bh30_w50_19 & '0' & '0' & '0' & '0' & heap_bh30_w45_18 & '0' & '0' & heap_bh30_w42_18 & '0' & '0' & heap_bh30_w39_18 & '0' & '0' & '0' & heap_bh30_w35_15 & heap_bh30_w34_17 & '0' & '0' & heap_bh30_w31_16 & '0' & '0' & heap_bh30_w28_16 & '0' & '0' & '0' & '0' & heap_bh30_w23_13 & '0' & '0' & heap_bh30_w20_12 & '0' & '0' & '0' & '0' & '0' & '0' & '0' & heap_bh30_w12_10 & '0' & '0' & '0' & '0' & heap_bh30_w7_7 & heap_bh30_w6_7 & heap_bh30_w5_6 & heap_bh30_w4_5 & '0' & '0' & heap_bh30_w1_1 & heap_bh30_w0_1;
   finalAdderCin_bh30 <= '0';
      Adder_final30_0: IntAdder_181_f400_uid1117
      port map ( Cin => finalAdderCin_bh30,
                 R => finalAdderOut_bh30,
                 X => finalAdderIn0_bh30,
                 Y => finalAdderIn1_bh30);
   -- concatenate all the compressed chunks
   CompressionResult30 <= finalAdderOut_bh30;
   -- End of code generated by BitHeap::generateCompressorVHDL
   R <= CompressionResult30(179 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                  RightShifter_189_by_max_100_comb_uid1127
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2011)
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity RightShifter_189_by_max_100_comb_uid1127 is
   port ( X : in  std_logic_vector(188 downto 0);
          S : in  std_logic_vector(6 downto 0);
          R : out  std_logic_vector(288 downto 0)   );
end entity;

architecture arch of RightShifter_189_by_max_100_comb_uid1127 is
signal level0 :  std_logic_vector(188 downto 0);
signal ps :  std_logic_vector(6 downto 0);
signal level1 :  std_logic_vector(189 downto 0);
signal level2 :  std_logic_vector(191 downto 0);
signal level3 :  std_logic_vector(195 downto 0);
signal level4 :  std_logic_vector(203 downto 0);
signal level5 :  std_logic_vector(219 downto 0);
signal level6 :  std_logic_vector(251 downto 0);
signal level7 :  std_logic_vector(315 downto 0);
begin
   level0<= X;
   ps<= S;
   level1<=  (0 downto 0 => '0') & level0 when ps(0) = '1' else    level0 & (0 downto 0 => '0');
   level2<=  (1 downto 0 => '0') & level1 when ps(1) = '1' else    level1 & (1 downto 0 => '0');
   level3<=  (3 downto 0 => '0') & level2 when ps(2) = '1' else    level2 & (3 downto 0 => '0');
   level4<=  (7 downto 0 => '0') & level3 when ps(3) = '1' else    level3 & (7 downto 0 => '0');
   level5<=  (15 downto 0 => '0') & level4 when ps(4) = '1' else    level4 & (15 downto 0 => '0');
   level6<=  (31 downto 0 => '0') & level5 when ps(5) = '1' else    level5 & (31 downto 0 => '0');
   level7<=  (63 downto 0 => '0') & level6 when ps(6) = '1' else    level6 & (63 downto 0 => '0');
   R <= level7(315 downto 27);
end architecture;

--------------------------------------------------------------------------------
--                         PositMult_100_8_comb_uid2
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Raul Murillo, 2019
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity PositMult_100_8_comb_uid2 is
   port ( InputA : in  std_logic_vector(99 downto 0);
          InputB : in  std_logic_vector(99 downto 0);
          Output : out  std_logic_vector(99 downto 0)   );
end entity;

architecture arch of PositMult_100_8_comb_uid2 is
   component PositDecoder_100_8_comb_uid4 is
      port ( Input : in  std_logic_vector(99 downto 0);
             Sign : out  std_logic;
             Reg : out  std_logic_vector(7 downto 0);
             Exp : out  std_logic_vector(7 downto 0);
             Frac : out  std_logic_vector(89 downto 0);
             z : out  std_logic;
             inf : out  std_logic   );
   end component;

   component PositDecoder_100_8_comb_uid16 is
      port ( Input : in  std_logic_vector(99 downto 0);
             Sign : out  std_logic;
             Reg : out  std_logic_vector(7 downto 0);
             Exp : out  std_logic_vector(7 downto 0);
             Frac : out  std_logic_vector(89 downto 0);
             z : out  std_logic;
             inf : out  std_logic   );
   end component;

   component IntMultiplier_UsingDSP_90_90_180_unsigned_comb_uid28 is
      port ( X : in  std_logic_vector(89 downto 0);
             Y : in  std_logic_vector(89 downto 0);
             R : out  std_logic_vector(179 downto 0)   );
   end component;

   component RightShifter_189_by_max_100_comb_uid1127 is
      port ( X : in  std_logic_vector(188 downto 0);
             S : in  std_logic_vector(6 downto 0);
             R : out  std_logic_vector(288 downto 0)   );
   end component;

signal sign_A :  std_logic;
signal reg_A :  std_logic_vector(7 downto 0);
signal exp_A :  std_logic_vector(7 downto 0);
signal frac_A :  std_logic_vector(89 downto 0);
signal z_A :  std_logic;
signal inf_A :  std_logic;
signal sign_B :  std_logic;
signal reg_B :  std_logic_vector(7 downto 0);
signal exp_B :  std_logic_vector(7 downto 0);
signal frac_B :  std_logic_vector(89 downto 0);
signal z_B :  std_logic;
signal inf_B :  std_logic;
signal sf_A :  std_logic_vector(15 downto 0);
signal sf_B :  std_logic_vector(15 downto 0);
signal sign :  std_logic;
signal z :  std_logic;
signal inf :  std_logic;
signal frac_mult :  std_logic_vector(179 downto 0);
signal ovf_m :  std_logic;
signal normFrac :  std_logic_vector(180 downto 0);
signal sf_mult :  std_logic_vector(16 downto 0);
signal sf_sign :  std_logic;
signal nzero :  std_logic;
signal ExpBits :  std_logic_vector(7 downto 0);
signal RegimeAns_tmp :  std_logic_vector(6 downto 0);
signal RegimeAns :  std_logic_vector(6 downto 0);
signal ovf_reg :  std_logic;
signal FinalRegime :  std_logic_vector(6 downto 0);
signal ovf_regF :  std_logic;
signal FinalExp :  std_logic_vector(7 downto 0);
signal tmp1 :  std_logic_vector(188 downto 0);
signal tmp2 :  std_logic_vector(188 downto 0);
signal shift_neg :  std_logic_vector(6 downto 0);
signal shift_pos :  std_logic_vector(6 downto 0);
signal shifter_in :  std_logic_vector(188 downto 0);
signal shifter_S :  std_logic_vector(6 downto 0);
signal shifter_out :  std_logic_vector(288 downto 0);
signal tmp_ans :  std_logic_vector(98 downto 0);
signal LSB :  std_logic;
signal G :  std_logic;
signal R :  std_logic;
signal S :  std_logic;
signal round :  std_logic;
begin
------------------------------- Data Extraction -------------------------------
   decoderA: PositDecoder_100_8_comb_uid4
      port map ( Exp => exp_A,
                 Frac => frac_A,
                 Input => InputA,
                 Reg => reg_A,
                 Sign => sign_A,
                 inf => inf_A,
                 z => z_A);
   decoderB: PositDecoder_100_8_comb_uid16
      port map ( Exp => exp_B,
                 Frac => frac_B,
                 Input => InputB,
                 Reg => reg_B,
                 Sign => sign_B,
                 inf => inf_B,
                 z => z_B);
   -- Gather scale factors
   sf_A <= reg_A & exp_A;
   sf_B <= reg_B & exp_B;
---------------------- Sign and Special Cases Computation ----------------------
   sign <= sign_A XOR sign_B;
   z <= z_A OR z_B;
   inf <= inf_A OR inf_B;
--------------- Multiply the fractions, add the exponent values ---------------
   mult: IntMultiplier_UsingDSP_90_90_180_unsigned_comb_uid28
      port map ( R => frac_mult,
                 X => frac_A,
                 Y => frac_B);
   -- Adjust for overflow
   ovf_m <= frac_mult(frac_mult'high);
   normFrac <= frac_mult & '0' when ovf_m = '0' else '0' & frac_mult;
   sf_mult <= (sf_A(sf_A'high) & sf_A) + (sf_B(sf_B'high) & sf_B) + ovf_m;
   sf_sign <= sf_mult(sf_mult'high);
---------------------- Compute Regime and Exponent value ----------------------
   nzero <= '0' when frac_mult = 0 else '1';
   -- Unpack scaling factors
   ExpBits <= sf_mult(7 downto 0);
   RegimeAns_tmp <= sf_mult(14 downto 8);
   -- Get Regime's absolute value
   RegimeAns <= (NOT RegimeAns_tmp)+1 when sf_sign = '1' else RegimeAns_tmp;
   -- Check for Regime overflow
   ovf_reg <= RegimeAns(RegimeAns'high);
   FinalRegime <= '0' & "111111" when ovf_reg = '1' else RegimeAns;
   ovf_regF <= '1' when FinalRegime = ('0' & "111111") else '0';
   FinalExp <= "00000000" when ((ovf_reg = '1') OR (ovf_regF = '1') OR (nzero='0')) else ExpBits;
------------------------------- Packing Stage 1 -------------------------------
   tmp1 <= nzero & '0' & FinalExp & normFrac(178 downto 0);
   tmp2 <= '0' & nzero & FinalExp & normFrac(178 downto 0);
   shift_neg <= FinalRegime - 2 when (ovf_regF = '1') else FinalRegime - 1;
   shift_pos <= FinalRegime - 1 when (ovf_regF = '1') else FinalRegime;
   shifter_in <= tmp2 when sf_sign = '1' else tmp1;
   shifter_S <= shift_neg when sf_sign = '1' else shift_pos;
   RightShifterComponent: RightShifter_189_by_max_100_comb_uid1127
      port map ( R => shifter_out,
                 S => shifter_S,
                 X => shifter_in);
   tmp_ans <= shifter_out(288 downto 190);
--------------------- Packing Stage 2 - Unbiased Rounding ---------------------
   LSB <= shifter_out(190);
   G <= shifter_out(189);
   R <= shifter_out(188);
   S <= '0' when shifter_out(187 downto 0) = 0 else '1';
   round <= G AND (LSB OR R OR S) when NOT((ovf_reg OR ovf_regF) = '1') else '0';
   Output <= '1' & "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" when inf = '1' else "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000" when z = '1' else '0' & (tmp_ans + round) when sign = '0' else NOT('0' & (tmp_ans + round))+1;
end architecture;


LIBRARY ieee; 
LIBRARY ieee_proposed; 
USE ieee.std_logic_1164.all; 
USE ieee.std_logic_arith.all; 
USE ieee.std_logic_unsigned.all; 
USE ieee.std_logic_textio.all; 
 
LIBRARY std; 
USE std.textio.all; 
USE ieee_proposed.fixed_pkg.all; 
USE ieee_proposed.fixed_float_types.all; 
USE ieee_proposed.float_pkg.all; 
ENTITY PCSystem_22 IS
    GENERIC (MantissaBits :INTEGER := 15 ; ExponentBits :INTEGER := 7 ; NumberOfBits :INTEGER := 22 ; FlopocoBits :INTEGER := 2);
    PORT (
    clk:IN std_logic;
    rst:IN std_logic;
    enable:IN std_logic;
    v1:IN std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
    v2:IN std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
    v3:IN std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
    v4:IN std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
    v5:IN std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
    v6:IN std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
    v7:IN std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
    v8:IN std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
    v9:IN std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
    v10:IN std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
    v11:IN std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
    v12:IN std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
    v13:IN std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
    v14:IN std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
    v15:IN std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
    v16:IN std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
    vb1:IN std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
    vb2:IN std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
    vb3:IN std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
    vb4:IN std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
    vb5:IN std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
    vb6:IN std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
    vb7:IN std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
    vb8:IN std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
    vb9:IN std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
    vb10:IN std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
    vb11:IN std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
    vb12:IN std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
    vb13:IN std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
    vb14:IN std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
    vb15:IN std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
    vb16:IN std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
    vout:OUT std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0)
);
END PCSystem_22;

ARCHITECTURE rtl of PCSystem_22 IS

        SIGNAL mb_D_FFMultiplier2_2293_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier2293_Output_2955 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF2293_2955MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF2293_2955MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF2293_2955MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF2293_2955MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR2293_2955Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR2293_2955Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier2_1146_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1146_Output_1477 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1146_1477MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1146_1477MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1146_1477MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1146_1477MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1146_1477Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1146_1477Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder3_Input1_661_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder661_Output_2954 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF661_2954AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF661_2954AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF661_2954AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF661_2954AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder3_Input2_661_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder3_Input1_330_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder330_Output_1476 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF330_1476AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF330_1476AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF330_1476AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF330_1476AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder3_Input2_330_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier4_2292_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier2292_Output_2953 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF2292_2953MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF2292_2953MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF2292_2953MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF2292_2953MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR2292_2953Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR2292_2953Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier4_1719_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1719_Output_2215 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1719_2215MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1719_2215MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1719_2215MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1719_2215MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1719_2215Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1719_2215Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier4_1145_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1145_Output_1475 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1145_1475MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1145_1475MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1145_1475MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1145_1475MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1145_1475Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1145_1475Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier4_572_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier572_Output_737 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF572_737MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF572_737MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF572_737MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF572_737MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR572_737Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR572_737Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder5_Input1_660_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder660_Output_2952 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF660_2952AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF660_2952AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF660_2952AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF660_2952AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder5_Input2_660_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder5_Input1_495_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder495_Output_2214 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF495_2214AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF495_2214AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF495_2214AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF495_2214AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder5_Input2_495_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder5_Input1_329_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder329_Output_1474 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF329_1474AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF329_1474AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF329_1474AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF329_1474AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder5_Input2_329_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder5_Input1_164_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder164_Output_736 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF164_736AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF164_736AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF164_736AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF164_736AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder5_Input2_164_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier6_Input1_2291_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier2291_Output_2951 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF2291_2951MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF2291_2951MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF2291_2951MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF2291_2951MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier6_Input2_2291_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier6_Input1_2005_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier2005_Output_2583 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF2005_2583MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF2005_2583MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF2005_2583MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF2005_2583MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier6_Input2_2005_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier6_Input1_1718_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1718_Output_2213 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1718_2213MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1718_2213MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1718_2213MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1718_2213MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier6_Input2_1718_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier6_Input1_1432_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1432_Output_1845 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1432_1845MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1432_1845MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1432_1845MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1432_1845MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier6_Input2_1432_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier6_Input1_1144_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1144_Output_1473 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1144_1473MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1144_1473MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1144_1473MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1144_1473MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier6_Input2_1144_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier6_Input1_858_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier858_Output_1105 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF858_1105MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF858_1105MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF858_1105MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF858_1105MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier6_Input2_858_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier6_Input1_571_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier571_Output_735 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF571_735MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF571_735MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF571_735MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF571_735MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier6_Input2_571_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier6_Input1_285_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier285_Output_367 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF285_367MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF285_367MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF285_367MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF285_367MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier6_Input2_285_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder7_Input1_659_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder659_Output_2950 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF659_2950AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF659_2950AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF659_2950AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF659_2950AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder7_Input2_659_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier7_2110_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier2110_Output_2711 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF2110_2711MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF2110_2711MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF2110_2711MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF2110_2711MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR2110_2711Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR2110_2711Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder7_Input1_577_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder577_Output_2582 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF577_2582AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF577_2582AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF577_2582AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF577_2582AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder7_Input2_577_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier7_1824_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1824_Output_2343 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1824_2343MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1824_2343MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1824_2343MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1824_2343MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1824_2343Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1824_2343Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder7_Input1_494_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder494_Output_2212 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF494_2212AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF494_2212AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF494_2212AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF494_2212AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder7_Input2_494_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier7_1537_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1537_Output_1973 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1537_1973MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1537_1973MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1537_1973MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1537_1973MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1537_1973Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1537_1973Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder7_Input1_412_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder412_Output_1844 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF412_1844AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF412_1844AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF412_1844AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF412_1844AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder7_Input2_412_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier7_1251_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1251_Output_1605 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1251_1605MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1251_1605MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1251_1605MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1251_1605MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1251_1605Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1251_1605Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder7_Input1_328_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder328_Output_1472 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF328_1472AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF328_1472AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF328_1472AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF328_1472AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder7_Input2_328_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier7_963_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier963_Output_1233 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF963_1233MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF963_1233MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF963_1233MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF963_1233MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR963_1233Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR963_1233Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder7_Input1_246_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder246_Output_1104 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF246_1104AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF246_1104AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF246_1104AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF246_1104AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder7_Input2_246_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier7_677_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier677_Output_865 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF677_865MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF677_865MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF677_865MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF677_865MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR677_865Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR677_865Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder7_Input1_163_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder163_Output_734 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF163_734AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF163_734AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF163_734AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF163_734AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder7_Input2_163_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier7_390_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier390_Output_495 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF390_495MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF390_495MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF390_495MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF390_495MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR390_495Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR390_495Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder7_Input1_81_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder81_Output_366 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF81_366AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF81_366AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF81_366AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF81_366AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder7_Input2_81_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier7_104_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier104_Output_127 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF104_127MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF104_127MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF104_127MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF104_127MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR104_127Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR104_127Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier8_2290_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier2290_Output_2949 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier2290WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier2290WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier2290WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF2290_2949MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF2290_2949MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR2290_2949Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier8_2200_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier2200_Output_2830 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier2200WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier2200WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier2200WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF2200_2830MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF2200_2830MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR2200_2830Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFAdder8_Input1_600_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder600_Output_2710 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF600_2710AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF600_2710AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF600_2710AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF600_2710AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder8_Input2_600_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier8_2004_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier2004_Output_2581 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier2004WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier2004WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier2004WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF2004_2581MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF2004_2581MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR2004_2581Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier8_1914_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1914_Output_2462 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier1914WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1914WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier1914WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1914_2462MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1914_2462MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1914_2462Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFAdder8_Input1_518_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder518_Output_2342 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF518_2342AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF518_2342AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF518_2342AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF518_2342AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder8_Input2_518_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier8_1717_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1717_Output_2211 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier1717WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1717WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier1717WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1717_2211MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1717_2211MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1717_2211Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier8_1627_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1627_Output_2092 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier1627WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1627WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier1627WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1627_2092MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1627_2092MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1627_2092Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFAdder8_Input1_435_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder435_Output_1972 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF435_1972AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF435_1972AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF435_1972AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF435_1972AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder8_Input2_435_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier8_1431_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1431_Output_1843 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier1431WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1431WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier1431WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1431_1843MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1431_1843MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1431_1843Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier8_1341_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1341_Output_1724 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier1341WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1341WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier1341WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1341_1724MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1341_1724MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1341_1724Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFAdder8_Input1_353_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder353_Output_1604 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF353_1604AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF353_1604AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF353_1604AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF353_1604AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder8_Input2_353_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier8_1143_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1143_Output_1471 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier1143WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1143WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier1143WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1143_1471MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1143_1471MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1143_1471Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier8_1053_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1053_Output_1352 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier1053WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1053WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier1053WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1053_1352MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1053_1352MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1053_1352Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFAdder8_Input1_269_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder269_Output_1232 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF269_1232AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF269_1232AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF269_1232AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF269_1232AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder8_Input2_269_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier8_857_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier857_Output_1103 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier857WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier857WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier857WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF857_1103MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF857_1103MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR857_1103Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier8_767_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier767_Output_984 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier767WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier767WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier767WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF767_984MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF767_984MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR767_984Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFAdder8_Input1_187_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder187_Output_864 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF187_864AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF187_864AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF187_864AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF187_864AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder8_Input2_187_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier8_570_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier570_Output_733 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier570WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier570WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier570WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF570_733MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF570_733MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR570_733Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier8_480_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier480_Output_614 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier480WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier480WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier480WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF480_614MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF480_614MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR480_614Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFAdder8_Input1_104_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder104_Output_494 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF104_494AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF104_494AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF104_494AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF104_494AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder8_Input2_104_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier8_284_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier284_Output_365 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier284WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier284WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier284WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF284_365MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF284_365MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR284_365Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier8_194_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier194_Output_246 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier194WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier194WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier194WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF194_246MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF194_246MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR194_246Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFAdder8_Input1_22_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder22_Output_126 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF22_126AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF22_126AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF22_126AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF22_126AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder8_Input2_22_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier9_2003_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier2003_Output_2580 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF2003_2580MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF2003_2580MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF2003_2580MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF2003_2580MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR2003_2580Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR2003_2580Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier9_1913_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1913_Output_2461 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1913_2461MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1913_2461MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1913_2461MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1913_2461MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1913_2461Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1913_2461Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier9_2109_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier2109_Output_2709 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier2109WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier2109WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier2109WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF2109_2709MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF2109_2709MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR2109_2709Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier9_2057_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier2057_Output_2646 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier2057WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier2057WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier2057WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF2057_2646MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF2057_2646MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR2057_2646Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier9_1823_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1823_Output_2341 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier1823WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1823WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier1823WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1823_2341MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1823_2341MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1823_2341Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier9_1771_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1771_Output_2278 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier1771WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1771WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier1771WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1771_2278MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1771_2278MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1771_2278Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier9_1430_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1430_Output_1842 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1430_1842MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1430_1842MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1430_1842MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1430_1842MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1430_1842Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1430_1842Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier9_1340_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1340_Output_1723 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1340_1723MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1340_1723MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1340_1723MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1340_1723MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1340_1723Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1340_1723Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier9_1536_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1536_Output_1971 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier1536WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1536WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier1536WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1536_1971MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1536_1971MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1536_1971Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier9_1484_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1484_Output_1908 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier1484WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1484WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier1484WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1484_1908MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1484_1908MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1484_1908Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier9_1250_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1250_Output_1603 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier1250WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1250WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier1250WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1250_1603MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1250_1603MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1250_1603Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier9_1198_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1198_Output_1540 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier1198WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1198WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier1198WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1198_1540MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1198_1540MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1198_1540Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier9_856_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier856_Output_1102 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF856_1102MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF856_1102MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF856_1102MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF856_1102MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR856_1102Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR856_1102Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier9_766_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier766_Output_983 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF766_983MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF766_983MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF766_983MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF766_983MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR766_983Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR766_983Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier9_962_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier962_Output_1231 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier962WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier962WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier962WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF962_1231MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF962_1231MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR962_1231Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier9_910_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier910_Output_1168 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier910WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier910WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier910WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF910_1168MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF910_1168MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR910_1168Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier9_676_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier676_Output_863 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier676WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier676WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier676WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF676_863MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF676_863MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR676_863Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier9_624_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier624_Output_800 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier624WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier624WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier624WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF624_800MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF624_800MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR624_800Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier9_283_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier283_Output_364 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF283_364MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF283_364MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF283_364MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF283_364MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR283_364Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR283_364Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier9_193_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier193_Output_245 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF193_245MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF193_245MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF193_245MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF193_245MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR193_245Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR193_245Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier9_389_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier389_Output_493 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier389WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier389WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier389WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF389_493MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF389_493MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR389_493Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier9_337_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier337_Output_430 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier337WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier337WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier337WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF337_430MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF337_430MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR337_430Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier9_103_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier103_Output_125 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier103WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier103WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier103WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF103_125MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF103_125MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR103_125Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier9_51_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier51_Output_62 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier51WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier51WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier51WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF51_62MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF51_62MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR51_62Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFAdder10_Input1_576_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder576_Output_2579 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF576_2579AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF576_2579AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF576_2579AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF576_2579AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder10_Input2_576_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder10_Input1_547_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder547_Output_2460 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF547_2460AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF547_2460AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF547_2460AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF547_2460AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder10_Input2_547_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier10_961_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier961_Output_1230 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF961_1230MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF961_1230MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF961_1230MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF961_1230MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR961_1230Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR961_1230Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier10_909_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier909_Output_1167 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF909_1167MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF909_1167MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF909_1167MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF909_1167MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR909_1167Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR909_1167Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier10_675_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier675_Output_862 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF675_862MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF675_862MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF675_862MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF675_862MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR675_862Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR675_862Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier10_623_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier623_Output_799 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF623_799MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF623_799MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF623_799MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF623_799MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR623_799Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR623_799Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder10_Input1_411_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder411_Output_1841 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF411_1841AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF411_1841AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF411_1841AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF411_1841AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder10_Input2_411_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder10_Input1_382_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder382_Output_1722 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF382_1722AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF382_1722AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF382_1722AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF382_1722AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder10_Input2_382_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier10_388_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier388_Output_492 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF388_492MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF388_492MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF388_492MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF388_492MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR388_492Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR388_492Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier10_336_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier336_Output_429 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF336_429MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF336_429MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF336_429MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF336_429MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR336_429Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR336_429Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier10_102_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier102_Output_124 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF102_124MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF102_124MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF102_124MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF102_124MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR102_124Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR102_124Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier10_50_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier50_Output_61 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF50_61MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF50_61MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF50_61MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF50_61MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR50_61Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR50_61Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder10_Input1_245_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder245_Output_1101 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF245_1101AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF245_1101AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF245_1101AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF245_1101AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder10_Input2_245_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder10_Input1_216_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder216_Output_982 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF216_982AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF216_982AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF216_982AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF216_982AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder10_Input2_216_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder10_Input1_80_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder80_Output_363 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF80_363AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF80_363AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF80_363AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF80_363AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder10_Input2_80_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder10_Input1_51_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder51_Output_244 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF51_244AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF51_244AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF51_244AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF51_244AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder10_Input2_51_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier11_Input1_2002_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier2002_Output_2578 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF2002_2578MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF2002_2578MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF2002_2578MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF2002_2578MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier11_Input2_2002_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier11_Input1_1958_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1958_Output_2520 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1958_2520MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1958_2520MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1958_2520MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1958_2520MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier11_Input2_1958_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier11_Input1_1912_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1912_Output_2459 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1912_2459MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1912_2459MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1912_2459MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1912_2459MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier11_Input2_1912_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier11_Input1_1868_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1868_Output_2401 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1868_2401MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1868_2401MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1868_2401MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1868_2401MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier11_Input2_1868_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder11_Input1_268_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder268_Output_1229 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF268_1229AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF268_1229AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF268_1229AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF268_1229AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder11_Input2_268_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder11_Input1_257_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder257_Output_1166 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF257_1166AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF257_1166AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF257_1166AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF257_1166AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder11_Input2_257_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder11_Input1_186_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder186_Output_861 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF186_861AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF186_861AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF186_861AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF186_861AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder11_Input2_186_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder11_Input1_175_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder175_Output_798 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF175_798AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF175_798AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF175_798AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF175_798AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder11_Input2_175_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier11_Input1_1429_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1429_Output_1840 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1429_1840MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1429_1840MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1429_1840MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1429_1840MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier11_Input2_1429_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier11_Input1_1385_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1385_Output_1782 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1385_1782MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1385_1782MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1385_1782MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1385_1782MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier11_Input2_1385_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier11_Input1_1339_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1339_Output_1721 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1339_1721MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1339_1721MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1339_1721MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1339_1721MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier11_Input2_1339_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier11_Input1_1295_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1295_Output_1663 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1295_1663MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1295_1663MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1295_1663MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1295_1663MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier11_Input2_1295_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder11_Input1_103_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder103_Output_491 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF103_491AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF103_491AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF103_491AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF103_491AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder11_Input2_103_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder11_Input1_92_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder92_Output_428 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF92_428AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF92_428AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF92_428AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF92_428AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder11_Input2_92_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder11_Input1_21_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder21_Output_123 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF21_123AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF21_123AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF21_123AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF21_123AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder11_Input2_21_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder11_Input1_10_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder10_Output_60 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF10_60AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF10_60AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF10_60AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF10_60AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder11_Input2_10_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier11_Input1_855_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier855_Output_1100 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF855_1100MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF855_1100MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF855_1100MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF855_1100MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier11_Input2_855_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier11_Input1_811_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier811_Output_1042 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF811_1042MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF811_1042MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF811_1042MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF811_1042MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier11_Input2_811_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier11_Input1_765_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier765_Output_981 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF765_981MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF765_981MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF765_981MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF765_981MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier11_Input2_765_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier11_Input1_721_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier721_Output_923 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF721_923MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF721_923MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF721_923MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF721_923MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier11_Input2_721_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier11_Input1_282_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier282_Output_362 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF282_362MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF282_362MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF282_362MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF282_362MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier11_Input2_282_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier11_Input1_238_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier238_Output_304 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF238_304MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF238_304MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF238_304MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF238_304MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier11_Input2_238_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier11_Input1_192_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier192_Output_243 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF192_243MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF192_243MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF192_243MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF192_243MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier11_Input2_192_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier11_Input1_148_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier148_Output_185 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF148_185MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF148_185MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF148_185MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF148_185MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier11_Input2_148_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder12_Input1_410_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder410_Output_1839 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF410_1839AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF410_1839AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF410_1839AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF410_1839AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder12_Input2_410_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier12_844_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier844_Output_1086 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF844_1086MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF844_1086MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF844_1086MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF844_1086MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR844_1086Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR844_1086Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder12_Input1_396_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder396_Output_1781 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF396_1781AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF396_1781AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF396_1781AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF396_1781AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder12_Input2_396_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier12_800_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier800_Output_1028 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF800_1028MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF800_1028MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF800_1028MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF800_1028MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR800_1028Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR800_1028Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder12_Input1_381_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder381_Output_1720 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF381_1720AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF381_1720AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF381_1720AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF381_1720AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder12_Input2_381_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier12_754_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier754_Output_967 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF754_967MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF754_967MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF754_967MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF754_967MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR754_967Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR754_967Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder12_Input1_367_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder367_Output_1662 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF367_1662AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF367_1662AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF367_1662AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF367_1662AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder12_Input2_367_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier12_710_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier710_Output_909 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF710_909MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF710_909MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF710_909MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF710_909MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR710_909Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR710_909Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier12_960_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier960_Output_1228 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier960WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier960WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier960WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF960_1228MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF960_1228MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR960_1228Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier12_935_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier935_Output_1198 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier935WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier935WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier935WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF935_1198MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF935_1198MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR935_1198Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier12_908_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier908_Output_1165 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier908WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier908WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier908WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF908_1165MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF908_1165MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR908_1165Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier12_883_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier883_Output_1135 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier883WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier883WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier883WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF883_1135MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF883_1135MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR883_1135Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier12_674_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier674_Output_860 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier674WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier674WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier674WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF674_860MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF674_860MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR674_860Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier12_649_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier649_Output_830 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier649WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier649WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier649WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF649_830MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF649_830MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR649_830Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier12_622_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier622_Output_797 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier622WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier622WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier622WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF622_797MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF622_797MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR622_797Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier12_597_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier597_Output_767 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier597WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier597WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier597WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF597_767MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF597_767MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR597_767Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier12_271_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier271_Output_348 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF271_348MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF271_348MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF271_348MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF271_348MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR271_348Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR271_348Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier12_227_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier227_Output_290 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF227_290MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF227_290MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF227_290MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF227_290MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR227_290Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR227_290Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier12_181_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier181_Output_229 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF181_229MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF181_229MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF181_229MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF181_229MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR181_229Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR181_229Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier12_137_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier137_Output_171 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF137_171MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF137_171MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF137_171MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF137_171MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR137_171Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR137_171Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier12_387_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier387_Output_490 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier387WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier387WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier387WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF387_490MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF387_490MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR387_490Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier12_362_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier362_Output_460 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier362WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier362WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier362WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF362_460MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF362_460MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR362_460Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier12_335_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier335_Output_427 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier335WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier335WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier335WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF335_427MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF335_427MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR335_427Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier12_310_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier310_Output_397 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier310WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier310WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier310WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF310_397MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF310_397MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR310_397Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier12_101_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier101_Output_122 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier101WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier101WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier101WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF101_122MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF101_122MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR101_122Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier12_76_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier76_Output_92 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier76WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier76WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier76WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF76_92MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF76_92MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR76_92Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier12_49_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier49_Output_59 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier49WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier49WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier49WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF49_59MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF49_59MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR49_59Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier12_24_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier24_Output_29 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier24WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier24WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier24WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF24_29MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF24_29MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR24_29Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFAdder12_Input1_79_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder79_Output_361 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF79_361AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF79_361AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF79_361AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF79_361AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder12_Input2_79_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder12_Input1_65_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder65_Output_303 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF65_303AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF65_303AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF65_303AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF65_303AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder12_Input2_65_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder12_Input1_50_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder50_Output_242 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF50_242AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF50_242AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF50_242AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF50_242AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder12_Input2_50_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder12_Input1_36_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder36_Output_184 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF36_184AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF36_184AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF36_184AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF36_184AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder12_Input2_36_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier13_1428_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1428_Output_1838 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier1428WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1428WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier1428WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1428_1838MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1428_1838MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1428_1838Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier13_1423_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1423_Output_1832 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier1423WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1423WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier1423WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1423_1832MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1423_1832MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1423_1832Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFAdder13_Input1_241_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder241_Output_1085 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF241_1085AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF241_1085AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF241_1085AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF241_1085AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder13_Input2_241_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier13_1384_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1384_Output_1780 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier1384WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1384WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier1384WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1384_1780MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1384_1780MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1384_1780Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier13_1379_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1379_Output_1774 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier1379WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1379WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier1379WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1379_1774MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1379_1774MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1379_1774Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFAdder13_Input1_227_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder227_Output_1027 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF227_1027AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF227_1027AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF227_1027AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF227_1027AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder13_Input2_227_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier13_1338_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1338_Output_1719 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier1338WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1338WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier1338WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1338_1719MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1338_1719MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1338_1719Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier13_1333_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1333_Output_1713 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier1333WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1333WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier1333WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1333_1713MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1333_1713MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1333_1713Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFAdder13_Input1_212_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder212_Output_966 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF212_966AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF212_966AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF212_966AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF212_966AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder13_Input2_212_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier13_1294_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1294_Output_1661 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier1294WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1294WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier1294WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1294_1661MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1294_1661MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1294_1661Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier13_1289_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1289_Output_1655 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier1289WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1289WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier1289WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1289_1655MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1289_1655MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1289_1655Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFAdder13_Input1_198_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder198_Output_908 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF198_908AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF198_908AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF198_908AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF198_908AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder13_Input2_198_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier13_Input1_673_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier673_Output_859 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF673_859MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF673_859MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF673_859MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF673_859MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier13_Input2_673_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier13_Input1_648_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier648_Output_829 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF648_829MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF648_829MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF648_829MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF648_829MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier13_Input2_648_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier13_Input1_621_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier621_Output_796 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF621_796MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF621_796MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF621_796MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF621_796MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier13_Input2_621_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier13_Input1_596_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier596_Output_766 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF596_766MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF596_766MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF596_766MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF596_766MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier13_Input2_596_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder13_Input1_76_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder76_Output_347 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF76_347AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF76_347AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF76_347AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF76_347AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder13_Input2_76_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder13_Input1_62_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder62_Output_289 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF62_289AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF62_289AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF62_289AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF62_289AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder13_Input2_62_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder13_Input1_47_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder47_Output_228 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF47_228AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF47_228AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF47_228AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF47_228AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder13_Input2_47_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder13_Input1_33_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder33_Output_170 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF33_170AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF33_170AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF33_170AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF33_170AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder13_Input2_33_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier13_Input1_100_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier100_Output_121 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF100_121MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF100_121MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF100_121MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF100_121MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier13_Input2_100_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier13_Input1_75_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier75_Output_91 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF75_91MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF75_91MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF75_91MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF75_91MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier13_Input2_75_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier13_Input1_48_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier48_Output_58 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF48_58MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF48_58MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF48_58MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF48_58MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier13_Input2_48_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier13_Input1_23_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier23_Output_28 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF23_28MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF23_28MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF23_28MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF23_28MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier13_Input2_23_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier13_281_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier281_Output_360 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier281WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier281WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier281WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF281_360MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF281_360MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR281_360Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier13_276_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier276_Output_354 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier276WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier276WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier276WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF276_354MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF276_354MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR276_354Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier13_237_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier237_Output_302 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier237WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier237WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier237WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF237_302MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF237_302MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR237_302Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier13_232_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier232_Output_296 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier232WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier232WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier232WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF232_296MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF232_296MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR232_296Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier13_191_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier191_Output_241 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier191WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier191WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier191WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF191_241MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF191_241MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR191_241Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier13_186_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier186_Output_235 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier186WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier186WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier186WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF186_235MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF186_235MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR186_235Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier13_147_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier147_Output_183 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier147WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier147WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier147WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF147_183MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF147_183MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR147_183Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier13_142_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier142_Output_177 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier142WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier142WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier142WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF142_177MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF142_177MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR142_177Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier14_1427_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1427_Output_1837 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier1427WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1427WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier1427WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1427_1837MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1427_1837MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1427_1837Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier14_1422_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1422_Output_1831 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier1422WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1422WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier1422WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1422_1831MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1422_1831MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1422_1831Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier14_843_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier843_Output_1084 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier843WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier843WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier843WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF843_1084MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF843_1084MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR843_1084Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier14_827_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier827_Output_1063 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier827WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier827WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier827WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF827_1063MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF827_1063MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR827_1063Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier14_1383_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1383_Output_1779 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier1383WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1383WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier1383WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1383_1779MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1383_1779MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1383_1779Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier14_1378_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1378_Output_1773 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier1378WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1378WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier1378WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1378_1773MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1378_1773MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1378_1773Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier14_799_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier799_Output_1026 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier799WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier799WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier799WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF799_1026MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF799_1026MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR799_1026Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier14_783_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier783_Output_1005 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier783WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier783WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier783WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF783_1005MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF783_1005MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR783_1005Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier14_1337_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1337_Output_1718 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier1337WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1337WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier1337WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1337_1718MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1337_1718MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1337_1718Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier14_1332_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1332_Output_1712 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier1332WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1332WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier1332WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1332_1712MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1332_1712MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1332_1712Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier14_753_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier753_Output_965 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier753WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier753WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier753WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF753_965MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF753_965MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR753_965Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier14_737_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier737_Output_944 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier737WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier737WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier737WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF737_944MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF737_944MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR737_944Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier14_1293_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1293_Output_1660 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier1293WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1293WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier1293WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1293_1660MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1293_1660MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1293_1660Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier14_1288_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1288_Output_1654 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier1288WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1288WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier1288WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1288_1654MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1288_1654MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1288_1654Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier14_709_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier709_Output_907 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier709WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier709WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier709WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF709_907MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF709_907MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR709_907Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier14_693_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier693_Output_886 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier693WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier693WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier693WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF693_886MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF693_886MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR693_886Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFAdder14_Input1_185_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder185_Output_858 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF185_858AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF185_858AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF185_858AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF185_858AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder14_Input2_185_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier25_Output_30 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier25WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier25WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier25WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF25_30MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF25_30MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR25_Input1_30Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR25_Input2_30Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR25_Input2_30Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder14_Input1_180_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder180_Output_828 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF180_828AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF180_828AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF180_828AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF180_828AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder14_Input2_180_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier0_Output_0 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier0WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier0WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier0WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF0_0MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF0_0MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR0_Input1_0Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR0_Input2_0Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR0_Input2_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder14_Input1_174_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder174_Output_795 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF174_795AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF174_795AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF174_795AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF174_795AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder14_Input2_174_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder14_Input1_169_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder169_Output_765 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF169_765AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF169_765AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF169_765AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF169_765AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder14_Input2_169_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier14_270_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier270_Output_346 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier270WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier270WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier270WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF270_346MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF270_346MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR270_346Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier14_254_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier254_Output_325 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier254WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier254WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier254WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF254_325MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF254_325MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR254_325Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier14_226_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier226_Output_288 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier226WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier226WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier226WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF226_288MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF226_288MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR226_288Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier14_210_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier210_Output_267 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier210WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier210WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier210WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF210_267MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF210_267MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR210_267Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier14_180_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier180_Output_227 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier180WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier180WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier180WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF180_227MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF180_227MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR180_227Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier14_164_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier164_Output_206 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier164WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier164WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier164WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF164_206MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF164_206MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR164_206Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier14_136_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier136_Output_169 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier136WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier136WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier136WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF136_169MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF136_169MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR136_169Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier14_120_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier120_Output_148 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier120WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier120WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier120WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF120_148MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF120_148MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR120_148Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFAdder14_Input1_20_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder20_Output_120 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF20_120AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF20_120AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF20_120AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF20_120AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder14_Input2_20_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder14_Input1_15_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder15_Output_90 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF15_90AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF15_90AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF15_90AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF15_90AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder14_Input2_15_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder14_Input1_9_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder9_Output_57 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF9_57AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF9_57AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF9_57AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF9_57AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder14_Input2_9_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder14_Input1_4_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder4_Output_27 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF4_27AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF4_27AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF4_27AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF4_27AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder14_Input2_4_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier14_280_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier280_Output_359 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier280WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier280WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier280WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF280_359MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF280_359MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR280_359Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier14_275_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier275_Output_353 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier275WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier275WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier275WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF275_353MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF275_353MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR275_353Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier14_236_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier236_Output_301 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier236WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier236WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier236WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF236_301MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF236_301MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR236_301Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier14_231_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier231_Output_295 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier231WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier231WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier231WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF231_295MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF231_295MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR231_295Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier14_190_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier190_Output_240 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier190WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier190WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier190WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF190_240MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF190_240MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR190_240Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier14_185_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier185_Output_234 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier185WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier185WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier185WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF185_234MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF185_234MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR185_234Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier14_146_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier146_Output_182 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier146WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier146WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier146WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF146_182MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF146_182MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR146_182Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier14_141_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier141_Output_176 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier141WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier141WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier141WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF141_176MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF141_176MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR141_176Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier15_1336_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1336_Output_1717 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1336_1717MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1336_1717MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1336_1717MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1336_1717MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1336_1717Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1336_1717Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier15_1331_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1331_Output_1711 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1331_1711MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1331_1711MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1331_1711MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1331_1711MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1331_1711Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1331_1711Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier15_798_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier798_Output_1025 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF798_1025MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF798_1025MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF798_1025MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF798_1025MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR798_1025Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR798_1025Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier15_782_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier782_Output_1004 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF782_1004MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF782_1004MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF782_1004MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF782_1004MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR782_1004Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR782_1004Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier15_1292_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1292_Output_1659 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1292_1659MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1292_1659MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1292_1659MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1292_1659MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1292_1659Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1292_1659Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier15_1287_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1287_Output_1653 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1287_1653MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1287_1653MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1287_1653MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1287_1653MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1287_1653Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1287_1653Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier15_708_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier708_Output_906 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF708_906MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF708_906MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF708_906MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF708_906MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR708_906Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR708_906Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier15_692_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier692_Output_885 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF692_885MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF692_885MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF692_885MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF692_885MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR692_885Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR692_885Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier15_672_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier672_Output_857 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier672WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier672WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier672WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF672_857MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF672_857MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR672_857Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier15_661_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier661_Output_844 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier661WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier661WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier661WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF661_844MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF661_844MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR661_844Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier15_647_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier647_Output_827 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier647WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier647WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier647WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF647_827MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF647_827MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR647_827Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier15_636_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier636_Output_814 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier636WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier636WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier636WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF636_814MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF636_814MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR636_814Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier15_620_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier620_Output_794 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier620WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier620WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier620WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF620_794MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF620_794MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR620_794Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier15_609_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier609_Output_781 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier609WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier609WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier609WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF609_781MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF609_781MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR609_781Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier15_595_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier595_Output_764 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier595WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier595WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier595WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF595_764MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF595_764MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR595_764Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier15_584_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier584_Output_751 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier584WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier584WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier584WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF584_751MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF584_751MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR584_751Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier15_225_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier225_Output_287 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF225_287MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF225_287MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF225_287MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF225_287MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR225_287Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR225_287Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier15_209_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier209_Output_266 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF209_266MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF209_266MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF209_266MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF209_266MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR209_266Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR209_266Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier15_135_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier135_Output_168 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF135_168MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF135_168MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF135_168MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF135_168MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR135_168Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR135_168Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier15_119_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier119_Output_147 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF119_147MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF119_147MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF119_147MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF119_147MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR119_147Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR119_147Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier15_99_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier99_Output_119 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier99WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier99WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier99WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF99_119MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF99_119MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR99_119Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier15_88_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier88_Output_106 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier88WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier88WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier88WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF88_106MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF88_106MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR88_106Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier15_74_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier74_Output_89 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier74WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier74WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier74WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF74_89MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF74_89MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR74_89Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier15_63_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier63_Output_76 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier63WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier63WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier63WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF63_76MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF63_76MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR63_76Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier15_47_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier47_Output_56 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier47WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier47WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier47WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF47_56MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF47_56MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR47_56Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier15_36_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier36_Output_43 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier36WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier36WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier36WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF36_43MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF36_43MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR36_43Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier15_22_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier22_Output_26 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier22WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier22WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier22WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF22_26MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF22_26MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR22_26Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier15_11_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier11_Output_13 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier11WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier11WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier11WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF11_13MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF11_13MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR11_13Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier15_189_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier189_Output_239 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF189_239MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF189_239MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF189_239MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF189_239MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR189_239Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR189_239Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier15_184_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier184_Output_233 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF184_233MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF184_233MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF184_233MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF184_233MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR184_233Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR184_233Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier15_145_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier145_Output_181 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF145_181MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF145_181MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF145_181MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF145_181MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR145_181Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR145_181Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier15_140_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier140_Output_175 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF140_175MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF140_175MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF140_175MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF140_175MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR140_175Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR140_175Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder16_Input1_380_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder380_Output_1716 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF380_1716AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF380_1716AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF380_1716AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF380_1716AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder16_Input2_380_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder16_Input1_379_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder379_Output_1710 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF379_1710AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF379_1710AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF379_1710AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF379_1710AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder16_Input2_379_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder16_Input1_226_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder226_Output_1024 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF226_1024AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF226_1024AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF226_1024AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF226_1024AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder16_Input2_226_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder16_Input1_221_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder221_Output_1003 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF221_1003AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF221_1003AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF221_1003AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF221_1003AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder16_Input2_221_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder16_Input1_366_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder366_Output_1658 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF366_1658AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF366_1658AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF366_1658AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF366_1658AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder16_Input2_366_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder16_Input1_365_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder365_Output_1652 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF365_1652AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF365_1652AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF365_1652AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF365_1652AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder16_Input2_365_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder16_Input1_197_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder197_Output_905 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF197_905AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF197_905AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF197_905AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF197_905AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder16_Input2_197_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder16_Input1_192_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder192_Output_884 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF192_884AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF192_884AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF192_884AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF192_884AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder16_Input2_192_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier16_Input1_98_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier98_Output_118 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF98_118MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF98_118MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF98_118MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF98_118MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier16_Input2_98_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier16_Input1_87_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier87_Output_105 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF87_105MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF87_105MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF87_105MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF87_105MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier16_Input2_87_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier16_Input1_73_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier73_Output_88 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF73_88MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF73_88MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF73_88MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF73_88MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier16_Input2_73_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier16_Input1_62_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier62_Output_75 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF62_75MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF62_75MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF62_75MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF62_75MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier16_Input2_62_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier16_Input1_46_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier46_Output_55 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF46_55MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF46_55MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF46_55MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF46_55MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier16_Input2_46_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier16_Input1_35_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier35_Output_42 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF35_42MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF35_42MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF35_42MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF35_42MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier16_Input2_35_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier16_Input1_21_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier21_Output_25 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF21_25MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF21_25MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF21_25MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF21_25MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier16_Input2_21_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier16_Input1_10_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier10_Output_12 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF10_12MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF10_12MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF10_12MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF10_12MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier16_Input2_10_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder16_Input1_61_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder61_Output_286 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF61_286AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF61_286AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF61_286AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF61_286AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder16_Input2_61_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder16_Input1_56_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder56_Output_265 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF56_265AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF56_265AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF56_265AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF56_265AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder16_Input2_56_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder16_Input1_32_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder32_Output_167 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF32_167AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF32_167AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF32_167AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF32_167AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder16_Input2_32_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder16_Input1_27_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder27_Output_146 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF27_146AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF27_146AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF27_146AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF27_146AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder16_Input2_27_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder16_Input1_49_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder49_Output_238 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF49_238AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF49_238AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF49_238AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF49_238AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder16_Input2_49_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder16_Input1_48_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder48_Output_232 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF48_232AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF48_232AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF48_232AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF48_232AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder16_Input2_48_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder16_Input1_35_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder35_Output_180 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF35_180AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF35_180AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF35_180AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF35_180AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder16_Input2_35_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder16_Input1_34_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder34_Output_174 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF34_174AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF34_174AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF34_174AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF34_174AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder16_Input2_34_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1335_Output_1715 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier1335WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1335WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier1335WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1335_1715MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1335_1715MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1335_Input1_1715Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR1335_Input2_1715Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1335_Input2_1715Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1334_Output_1714 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier1334WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1334WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier1334WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1334_1714MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1334_1714MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1334_Input1_1714Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR1334_Input2_1714Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1334_Input2_1714Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1330_Output_1709 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier1330WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1330WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier1330WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1330_1709MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1330_1709MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1330_Input1_1709Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR1330_Input2_1709Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1330_Input2_1709Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1329_Output_1708 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier1329WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1329WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier1329WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1329_1708MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1329_1708MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1329_Input1_1708Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR1329_Input2_1708Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1329_Input2_1708Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier17_Input1_797_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier797_Output_1023 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF797_1023MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF797_1023MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF797_1023MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF797_1023MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier17_Input2_797_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier17_Input1_790_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier790_Output_1014 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF790_1014MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF790_1014MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF790_1014MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF790_1014MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier17_Input2_790_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier17_Input1_781_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier781_Output_1002 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF781_1002MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF781_1002MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF781_1002MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF781_1002MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier17_Input2_781_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier17_Input1_774_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier774_Output_993 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF774_993MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF774_993MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF774_993MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF774_993MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier17_Input2_774_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1291_Output_1657 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier1291WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1291WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier1291WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1291_1657MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1291_1657MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1291_Input1_1657Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR1291_Input2_1657Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1291_Input2_1657Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1290_Output_1656 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier1290WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1290WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier1290WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1290_1656MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1290_1656MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1290_Input1_1656Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR1290_Input2_1656Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1290_Input2_1656Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1286_Output_1651 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier1286WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1286WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier1286WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1286_1651MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1286_1651MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1286_Input1_1651Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR1286_Input2_1651Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1286_Input2_1651Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1285_Output_1650 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier1285WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1285WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier1285WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1285_1650MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1285_1650MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1285_Input1_1650Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR1285_Input2_1650Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1285_Input2_1650Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier17_Input1_707_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier707_Output_904 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF707_904MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF707_904MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF707_904MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF707_904MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier17_Input2_707_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier17_Input1_700_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier700_Output_895 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF700_895MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF700_895MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF700_895MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF700_895MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier17_Input2_700_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier17_Input1_691_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier691_Output_883 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF691_883MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF691_883MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF691_883MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF691_883MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier17_Input2_691_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier17_Input1_684_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier684_Output_874 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF684_874MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF684_874MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF684_874MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF684_874MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier17_Input2_684_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder17_Input1_19_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder19_Output_117 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF19_117AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF19_117AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF19_117AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF19_117AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder17_Input2_19_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier17_91_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier91_Output_110 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF91_110MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF91_110MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF91_110MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF91_110MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR91_110Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR91_110Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder17_Input1_17_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder17_Output_104 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF17_104AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF17_104AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF17_104AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF17_104AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder17_Input2_17_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier17_80_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier80_Output_97 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF80_97MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF80_97MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF80_97MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF80_97MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR80_97Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR80_97Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder17_Input1_14_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder14_Output_87 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF14_87AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF14_87AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF14_87AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF14_87AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder17_Input2_14_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier17_66_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier66_Output_80 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF66_80MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF66_80MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF66_80MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF66_80MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR66_80Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR66_80Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder17_Input1_12_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder12_Output_74 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF12_74AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF12_74AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF12_74AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF12_74AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder17_Input2_12_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier17_55_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier55_Output_67 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF55_67MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF55_67MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF55_67MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF55_67MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR55_67Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR55_67Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder17_Input1_8_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder8_Output_54 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF8_54AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF8_54AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF8_54AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF8_54AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder17_Input2_8_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier17_39_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier39_Output_47 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF39_47MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF39_47MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF39_47MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF39_47MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR39_47Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR39_47Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder17_Input1_6_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder6_Output_41 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF6_41AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF6_41AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF6_41AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF6_41AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder17_Input2_6_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier17_28_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier28_Output_34 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF28_34MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF28_34MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF28_34MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF28_34MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR28_34Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR28_34Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder17_Input1_3_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder3_Output_24 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF3_24AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF3_24AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF3_24AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF3_24AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder17_Input2_3_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier17_14_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier14_Output_17 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF14_17MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF14_17MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF14_17MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF14_17MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR14_17Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR14_17Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder17_Input1_1_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder1_Output_11 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1_11AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1_11AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1_11AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1_11AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder17_Input2_1_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier17_3_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier3_Output_4 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF3_4MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF3_4MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF3_4MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF3_4MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR3_4Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR3_4Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier17_Input1_224_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier224_Output_285 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF224_285MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF224_285MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF224_285MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF224_285MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier17_Input2_224_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier17_Input1_217_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier217_Output_276 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF217_276MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF217_276MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF217_276MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF217_276MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier17_Input2_217_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier17_Input1_208_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier208_Output_264 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF208_264MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF208_264MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF208_264MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF208_264MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier17_Input2_208_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier17_Input1_201_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier201_Output_255 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF201_255MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF201_255MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF201_255MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF201_255MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier17_Input2_201_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier17_Input1_134_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier134_Output_166 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF134_166MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF134_166MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF134_166MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF134_166MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier17_Input2_134_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier17_Input1_127_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier127_Output_157 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF127_157MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF127_157MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF127_157MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF127_157MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier17_Input2_127_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier17_Input1_118_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier118_Output_145 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF118_145MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF118_145MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF118_145MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF118_145MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier17_Input2_118_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier17_Input1_111_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier111_Output_136 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF111_136MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF111_136MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF111_136MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF111_136MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier17_Input2_111_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier188_Output_237 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier188WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier188WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier188WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF188_237MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF188_237MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR188_Input1_237Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR188_Input2_237Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR188_Input2_237Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier187_Output_236 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier187WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier187WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier187WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF187_236MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF187_236MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR187_Input1_236Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR187_Input2_236Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR187_Input2_236Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier183_Output_231 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier183WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier183WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier183WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF183_231MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF183_231MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR183_Input1_231Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR183_Input2_231Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR183_Input2_231Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier182_Output_230 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier182WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier182WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier182WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF182_230MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF182_230MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR182_Input1_230Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR182_Input2_230Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR182_Input2_230Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier144_Output_179 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier144WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier144WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier144WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF144_179MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF144_179MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR144_Input1_179Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR144_Input2_179Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR144_Input2_179Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier143_Output_178 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier143WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier143WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier143WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF143_178MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF143_178MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR143_Input1_178Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR143_Input2_178Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR143_Input2_178Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier139_Output_173 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier139WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier139WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier139WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF139_173MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF139_173MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR139_Input1_173Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR139_Input2_173Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR139_Input2_173Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier138_Output_172 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier138WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier138WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier138WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF138_172MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF138_172MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR138_Input1_172Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR138_Input2_172Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR138_Input2_172Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder18_Input1_60_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder60_Output_284 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF60_284AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF60_284AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF60_284AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF60_284AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder18_Input2_60_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier18_704_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier704_Output_900 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier704WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier704WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier704WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF704_900MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF704_900MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR704_900Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFAdder18_Input1_58_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder58_Output_275 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF58_275AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF58_275AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF58_275AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF58_275AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder18_Input2_58_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier18_697_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier697_Output_891 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier697WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier697WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier697WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF697_891MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF697_891MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR697_891Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFAdder18_Input1_55_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder55_Output_263 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF55_263AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF55_263AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF55_263AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF55_263AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder18_Input2_55_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier18_688_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier688_Output_879 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier688WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier688WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier688WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF688_879MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF688_879MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR688_879Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFAdder18_Input1_53_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder53_Output_254 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF53_254AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF53_254AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF53_254AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF53_254AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder18_Input2_53_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier18_681_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier681_Output_870 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier681WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier681WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier681WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF681_870MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF681_870MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR681_870Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFAdder18_Input1_31_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder31_Output_165 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF31_165AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF31_165AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF31_165AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF31_165AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder18_Input2_31_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder18_Input1_29_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder29_Output_156 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF29_156AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF29_156AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF29_156AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF29_156AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder18_Input2_29_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder18_Input1_26_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder26_Output_144 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF26_144AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF26_144AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF26_144AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF26_144AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder18_Input2_26_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder18_Input1_24_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder24_Output_135 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF24_135AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF24_135AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF24_135AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF24_135AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder18_Input2_24_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier18_97_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier97_Output_116 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier97WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier97WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier97WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF97_116MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF97_116MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR97_116Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier18_94_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier94_Output_113 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier94WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier94WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier94WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF94_113MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF94_113MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR94_113Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFAdder18_Input1_18_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder18_Output_109 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF18_109AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF18_109AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF18_109AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF18_109AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder18_Input2_18_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier18_86_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier86_Output_103 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier86WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier86WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier86WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF86_103MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF86_103MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR86_103Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier18_83_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier83_Output_100 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier83WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier83WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier83WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF83_100MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF83_100MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR83_100Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFAdder18_Input1_16_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder16_Output_96 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF16_96AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF16_96AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF16_96AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF16_96AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder18_Input2_16_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier18_72_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier72_Output_86 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier72WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier72WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier72WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF72_86MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF72_86MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR72_86Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier18_69_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier69_Output_83 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier69WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier69WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier69WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF69_83MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF69_83MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR69_83Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFAdder18_Input1_13_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder13_Output_79 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF13_79AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF13_79AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF13_79AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF13_79AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder18_Input2_13_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier18_61_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier61_Output_73 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier61WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier61WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier61WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF61_73MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF61_73MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR61_73Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier18_58_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier58_Output_70 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier58WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier58WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier58WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF58_70MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF58_70MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR58_70Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFAdder18_Input1_11_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder11_Output_66 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF11_66AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF11_66AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF11_66AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF11_66AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder18_Input2_11_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier18_45_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier45_Output_53 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier45WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier45WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier45WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF45_53MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF45_53MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR45_53Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier18_42_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier42_Output_50 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier42WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier42WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier42WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF42_50MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF42_50MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR42_50Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFAdder18_Input1_7_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder7_Output_46 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF7_46AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF7_46AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF7_46AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF7_46AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder18_Input2_7_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier18_34_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier34_Output_40 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier34WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier34WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier34WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF34_40MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF34_40MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR34_40Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier18_31_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier31_Output_37 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier31WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier31WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier31WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF31_37MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF31_37MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR31_37Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFAdder18_Input1_5_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder5_Output_33 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF5_33AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF5_33AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF5_33AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF5_33AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder18_Input2_5_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier18_20_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier20_Output_23 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier20WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier20WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier20WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF20_23MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF20_23MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR20_23Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier18_17_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier17_Output_20 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier17WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier17WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier17WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF17_20MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF17_20MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR17_20Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFAdder18_Input1_2_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder2_Output_16 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF2_16AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF2_16AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF2_16AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF2_16AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder18_Input2_2_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier18_9_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier9_Output_10 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier9WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier9WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier9WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF9_10MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF9_10MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR9_10Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier18_6_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier6_Output_7 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier6WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier6WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier6WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF6_7MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF6_7MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR6_7Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFAdder18_Input1_0_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder0_Output_3 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF0_3AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF0_3AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF0_3AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF0_3AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder18_Input2_0_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier18_131_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier131_Output_162 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier131WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier131WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier131WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF131_162MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF131_162MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR131_162Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier18_124_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier124_Output_153 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier124WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier124WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier124WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF124_153MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF124_153MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR124_153Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier18_115_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier115_Output_141 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier115WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier115WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier115WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF115_141MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF115_141MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR115_141Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier18_108_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier108_Output_132 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier108WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier108WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier108WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF108_132MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF108_132MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR108_132Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL Multiplier223_Output_283 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier223WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier223WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier223WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF223_283MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF223_283MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR223_Input1_283Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR223_Input2_283Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR223_Input2_283Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier222_Output_282 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier222WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier222WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier222WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF222_282MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF222_282MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR222_Input1_282Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR222_Input2_282Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR222_Input2_282Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier19_703_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier703_Output_899 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF703_899MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF703_899MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF703_899MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF703_899MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR703_899Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR703_899Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier216_Output_274 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier216WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier216WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier216WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF216_274MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF216_274MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR216_Input1_274Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR216_Input2_274Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR216_Input2_274Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier215_Output_273 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier215WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier215WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier215WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF215_273MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF215_273MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR215_Input1_273Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR215_Input2_273Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR215_Input2_273Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier19_696_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier696_Output_890 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF696_890MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF696_890MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF696_890MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF696_890MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR696_890Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR696_890Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier207_Output_262 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier207WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier207WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier207WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF207_262MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF207_262MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR207_Input1_262Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR207_Input2_262Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR207_Input2_262Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier206_Output_261 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier206WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier206WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier206WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF206_261MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF206_261MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR206_Input1_261Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR206_Input2_261Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR206_Input2_261Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier19_687_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier687_Output_878 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF687_878MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF687_878MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF687_878MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF687_878MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR687_878Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR687_878Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier200_Output_253 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier200WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier200WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier200WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF200_253MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF200_253MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR200_Input1_253Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR200_Input2_253Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR200_Input2_253Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier199_Output_252 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier199WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier199WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier199WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF199_252MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF199_252MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR199_Input1_252Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR199_Input2_252Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR199_Input2_252Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier19_680_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier680_Output_869 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF680_869MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF680_869MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF680_869MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF680_869MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR680_869Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR680_869Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier133_Output_164 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier133WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier133WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier133WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF133_164MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF133_164MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR133_Input1_164Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR133_Input2_164Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR133_Input2_164Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier132_Output_163 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier132WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier132WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier132WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF132_163MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF132_163MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR132_Input1_163Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR132_Input2_163Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR132_Input2_163Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier126_Output_155 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier126WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier126WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier126WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF126_155MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF126_155MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR126_Input1_155Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR126_Input2_155Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR126_Input2_155Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier125_Output_154 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier125WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier125WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier125WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF125_154MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF125_154MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR125_Input1_154Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR125_Input2_154Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR125_Input2_154Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier117_Output_143 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier117WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier117WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier117WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF117_143MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF117_143MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR117_Input1_143Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR117_Input2_143Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR117_Input2_143Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier116_Output_142 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier116WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier116WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier116WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF116_142MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF116_142MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR116_Input1_142Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR116_Input2_142Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR116_Input2_142Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier110_Output_134 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier110WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier110WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier110WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF110_134MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF110_134MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR110_Input1_134Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR110_Input2_134Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR110_Input2_134Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier109_Output_133 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier109WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier109WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier109WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF109_133MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF109_133MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR109_Input1_133Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR109_Input2_133Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR109_Input2_133Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier19_44_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier44_Output_52 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier44WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier44WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier44WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF44_52MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF44_52MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR44_52Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier19_41_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier41_Output_49 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier41WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier41WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier41WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF41_49MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF41_49MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR41_49Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL Multiplier90_Output_108 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier90WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier90WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier90WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF90_108MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF90_108MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR90_Input1_108Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR90_Input2_108Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR90_Input2_108Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier89_Output_107 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier89WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier89WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier89WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF89_107MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF89_107MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR89_Input1_107Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR89_Input2_107Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR89_Input2_107Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier19_33_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier33_Output_39 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier33WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier33WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier33WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF33_39MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF33_39MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR33_39Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier19_30_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier30_Output_36 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier30WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier30WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier30WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF30_36MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF30_36MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR30_36Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL Multiplier79_Output_95 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier79WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier79WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier79WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF79_95MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF79_95MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR79_Input1_95Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR79_Input2_95Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR79_Input2_95Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier78_Output_94 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier78WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier78WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier78WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF78_94MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF78_94MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR78_Input1_94Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR78_Input2_94Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR78_Input2_94Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier19_19_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier19_Output_22 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier19WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier19WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier19WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF19_22MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF19_22MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR19_22Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier19_16_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier16_Output_19 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier16WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier16WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier16WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF16_19MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF16_19MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR16_19Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL Multiplier65_Output_78 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier65WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier65WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier65WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF65_78MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF65_78MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR65_Input1_78Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR65_Input2_78Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR65_Input2_78Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier64_Output_77 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier64WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier64WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier64WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF64_77MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF64_77MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR64_Input1_77Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR64_Input2_77Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR64_Input2_77Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier19_8_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier8_Output_9 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier8WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier8WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier8WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF8_9MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF8_9MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR8_9Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier19_5_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier5_Output_6 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier5WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier5WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier5WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF5_6MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF5_6MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR5_6Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL Multiplier54_Output_65 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier54WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier54WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier54WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF54_65MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF54_65MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR54_Input1_65Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR54_Input2_65Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR54_Input2_65Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier53_Output_64 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier53WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier53WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier53WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF53_64MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF53_64MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR53_Input1_64Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR53_Input2_64Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR53_Input2_64Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier38_Output_45 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier38WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier38WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier38WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF38_45MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF38_45MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR38_Input1_45Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR38_Input2_45Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR38_Input2_45Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier37_Output_44 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier37WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier37WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier37WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF37_44MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF37_44MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR37_Input1_44Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR37_Input2_44Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR37_Input2_44Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier27_Output_32 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier27WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier27WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier27WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF27_32MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF27_32MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR27_Input1_32Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR27_Input2_32Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR27_Input2_32Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier26_Output_31 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier26WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier26WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier26WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF26_31MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF26_31MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR26_Input1_31Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR26_Input2_31Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR26_Input2_31Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier13_Output_15 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier13WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier13WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier13WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF13_15MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF13_15MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR13_Input1_15Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR13_Input2_15Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR13_Input2_15Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier12_Output_14 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier12WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier12WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier12WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF12_14MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF12_14MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR12_Input1_14Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR12_Input2_14Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR12_Input2_14Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier2_Output_2 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier2WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier2WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier2WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF2_2MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF2_2MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR2_Input1_2Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR2_Input2_2Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR2_Input2_2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1_Output_1 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier1WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier1WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1_1MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1_1MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1_Input1_1Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR1_Input2_1Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1_Input2_1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier19_130_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier130_Output_161 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF130_161MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF130_161MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF130_161MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF130_161MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR130_161Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR130_161Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier19_123_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier123_Output_152 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF123_152MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF123_152MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF123_152MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF123_152MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR123_152Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR123_152Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier19_114_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier114_Output_140 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF114_140MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF114_140MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF114_140MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF114_140MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR114_140Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR114_140Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier19_107_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier107_Output_131 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF107_131MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF107_131MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF107_131MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF107_131MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR107_131Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR107_131Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder20_Input1_195_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder195_Output_898 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF195_898AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF195_898AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF195_898AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF195_898AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder20_Input2_195_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder20_Input1_193_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder193_Output_889 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF193_889AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF193_889AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF193_889AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF193_889AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder20_Input2_193_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder20_Input1_190_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder190_Output_877 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF190_877AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF190_877AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF190_877AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF190_877AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder20_Input2_190_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder20_Input1_188_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder188_Output_868 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF188_868AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF188_868AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF188_868AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF188_868AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder20_Input2_188_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier32_Output_38 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier32WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier32WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier32WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF32_38MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF32_38MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR32_Input1_38Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR32_Input2_38Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR32_Input2_38Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier29_Output_35 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier29WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier29WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier29WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF29_35MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF29_35MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR29_Input1_35Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR29_Input2_35Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR29_Input2_35Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier7_Output_8 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier7WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier7WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier7WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF7_8MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF7_8MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR7_Input1_8Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR7_Input2_8Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR7_Input2_8Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier4_Output_5 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier4WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier4WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier4WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF4_5MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF4_5MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR4_Input1_5Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR4_Input2_5Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR4_Input2_5Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder20_Input1_30_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder30_Output_160 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF30_160AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF30_160AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF30_160AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF30_160AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder20_Input2_30_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder20_Input1_28_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder28_Output_151 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF28_151AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF28_151AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF28_151AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF28_151AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder20_Input2_28_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder20_Input1_25_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder25_Output_139 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF25_139AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF25_139AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF25_139AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF25_139AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder20_Input2_25_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder20_Input1_23_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder23_Output_130 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF23_130AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF23_130AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF23_130AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF23_130AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder20_Input2_23_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier702_Output_897 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier702WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier702WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier702WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF702_897MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF702_897MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR702_897Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier21_702_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier21_702_0Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier701_Output_896 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier701WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier701WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier701WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF701_896MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF701_896MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR701_896Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier21_701_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier21_701_0Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier695_Output_888 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier695WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier695WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier695WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF695_888MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF695_888MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR695_888Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier21_695_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier21_695_0Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier694_Output_887 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier694WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier694WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier694WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF694_887MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF694_887MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR694_887Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier21_694_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier21_694_0Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier686_Output_876 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier686WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier686WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier686WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF686_876MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF686_876MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR686_876Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier21_686_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier21_686_0Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier685_Output_875 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier685WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier685WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier685WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF685_875MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF685_875MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR685_875Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier21_685_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier21_685_0Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier679_Output_867 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier679WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier679WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier679WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF679_867MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF679_867MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR679_867Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier21_679_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier21_679_0Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier678_Output_866 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier678WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier678WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier678WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF678_866MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF678_866MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR678_866Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier21_678_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier21_678_0Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier129_Output_159 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier129WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier129WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier129WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF129_159MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF129_159MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR129_159Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier21_129_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier21_129_0Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier128_Output_158 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier128WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier128WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier128WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF128_158MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF128_158MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR128_158Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier21_128_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier21_128_0Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier122_Output_150 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier122WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier122WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier122WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF122_150MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF122_150MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR122_150Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier21_122_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier21_122_0Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier121_Output_149 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier121WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier121WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier121WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF121_149MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF121_149MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR121_149Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier21_121_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier21_121_0Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier113_Output_138 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier113WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier113WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier113WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF113_138MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF113_138MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR113_138Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier21_113_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier21_113_0Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier112_Output_137 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier112WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier112WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier112WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF112_137MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF112_137MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR112_137Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier21_112_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier21_112_0Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier106_Output_129 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier106WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier106WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier106WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF106_129MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF106_129MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR106_129Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier21_106_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier21_106_0Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier105_Output_128 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier105WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier105WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier105WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF105_128MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF105_128MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR105_128Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier21_105_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier21_105_0Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder1_Input1_662_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder662_Output_2956 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF662_2956AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF662_2956AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF662_2956AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF662_2956AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder1_Input2_662_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder1_Output_662_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier0Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.848299,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.895308,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.842608,exponentBits,mantissaBits-1));
        SIGNAL Multiplier4Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870697,exponentBits,mantissaBits-1));
        SIGNAL Multiplier5Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.945793,exponentBits,mantissaBits-1));
        SIGNAL Multiplier6Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.95487,exponentBits,mantissaBits-1));
        SIGNAL Multiplier7Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870404,exponentBits,mantissaBits-1));
        SIGNAL Multiplier8Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.780732,exponentBits,mantissaBits-1));
        SIGNAL Multiplier9Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.810846,exponentBits,mantissaBits-1));
        SIGNAL Multiplier11Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.991361,exponentBits,mantissaBits-1));
        SIGNAL Multiplier12Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.669241,exponentBits,mantissaBits-1));
        SIGNAL Multiplier13Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.97158,exponentBits,mantissaBits-1));
        SIGNAL Multiplier15Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870697,exponentBits,mantissaBits-1));
        SIGNAL Multiplier16Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.75369,exponentBits,mantissaBits-1));
        SIGNAL Multiplier17Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.77448,exponentBits,mantissaBits-1));
        SIGNAL Multiplier18Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870404,exponentBits,mantissaBits-1));
        SIGNAL Multiplier19Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.933776,exponentBits,mantissaBits-1));
        SIGNAL Multiplier20Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.660973,exponentBits,mantissaBits-1));
        SIGNAL Multiplier22Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870239,exponentBits,mantissaBits-1));
        SIGNAL Multiplier24Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.94472,exponentBits,mantissaBits-1));
        SIGNAL Multiplier25Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.890735,exponentBits,mantissaBits-1));
        SIGNAL Multiplier26Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.689002,exponentBits,mantissaBits-1));
        SIGNAL Multiplier27Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.966814,exponentBits,mantissaBits-1));
        SIGNAL Multiplier29Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.551341,exponentBits,mantissaBits-1));
        SIGNAL Multiplier30Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.795357,exponentBits,mantissaBits-1));
        SIGNAL Multiplier31Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.746308,exponentBits,mantissaBits-1));
        SIGNAL Multiplier32Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.989597,exponentBits,mantissaBits-1));
        SIGNAL Multiplier33Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.577708,exponentBits,mantissaBits-1));
        SIGNAL Multiplier34Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.618274,exponentBits,mantissaBits-1));
        SIGNAL Multiplier36Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.952809,exponentBits,mantissaBits-1));
        SIGNAL Multiplier37Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.495915,exponentBits,mantissaBits-1));
        SIGNAL Multiplier38Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.993928,exponentBits,mantissaBits-1));
        SIGNAL Multiplier40Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.551341,exponentBits,mantissaBits-1));
        SIGNAL Multiplier41Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.926235,exponentBits,mantissaBits-1));
        SIGNAL Multiplier42Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.616494,exponentBits,mantissaBits-1));
        SIGNAL Multiplier43Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.989597,exponentBits,mantissaBits-1));
        SIGNAL Multiplier44Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.986786,exponentBits,mantissaBits-1));
        SIGNAL Multiplier45Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.464416,exponentBits,mantissaBits-1));
        SIGNAL Multiplier47Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.770987,exponentBits,mantissaBits-1));
        SIGNAL Multiplier49Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.827729,exponentBits,mantissaBits-1));
        SIGNAL Multiplier51Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.986612,exponentBits,mantissaBits-1));
        SIGNAL Multiplier52Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.848299,exponentBits,mantissaBits-1));
        SIGNAL Multiplier53Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.562709,exponentBits,mantissaBits-1));
        SIGNAL Multiplier54Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.988453,exponentBits,mantissaBits-1));
        SIGNAL Multiplier56Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870697,exponentBits,mantissaBits-1));
        SIGNAL Multiplier57Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.945793,exponentBits,mantissaBits-1));
        SIGNAL Multiplier58Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.729204,exponentBits,mantissaBits-1));
        SIGNAL Multiplier59Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870404,exponentBits,mantissaBits-1));
        SIGNAL Multiplier60Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.780732,exponentBits,mantissaBits-1));
        SIGNAL Multiplier61Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.917308,exponentBits,mantissaBits-1));
        SIGNAL Multiplier63Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.979033,exponentBits,mantissaBits-1));
        SIGNAL Multiplier64Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.453222,exponentBits,mantissaBits-1));
        SIGNAL Multiplier65Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.996146,exponentBits,mantissaBits-1));
        SIGNAL Multiplier67Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870697,exponentBits,mantissaBits-1));
        SIGNAL Multiplier68Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.75369,exponentBits,mantissaBits-1));
        SIGNAL Multiplier69Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.936763,exponentBits,mantissaBits-1));
        SIGNAL Multiplier70Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870404,exponentBits,mantissaBits-1));
        SIGNAL Multiplier71Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.933776,exponentBits,mantissaBits-1));
        SIGNAL Multiplier72Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.973389,exponentBits,mantissaBits-1));
        SIGNAL Multiplier74Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.818419,exponentBits,mantissaBits-1));
        SIGNAL Multiplier76Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.766253,exponentBits,mantissaBits-1));
        SIGNAL Multiplier77Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.890735,exponentBits,mantissaBits-1));
        SIGNAL Multiplier78Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.382644,exponentBits,mantissaBits-1));
        SIGNAL Multiplier79Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.998354,exponentBits,mantissaBits-1));
        SIGNAL Multiplier81Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.551341,exponentBits,mantissaBits-1));
        SIGNAL Multiplier82Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.795357,exponentBits,mantissaBits-1));
        SIGNAL Multiplier83Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.948695,exponentBits,mantissaBits-1));
        SIGNAL Multiplier84Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.989597,exponentBits,mantissaBits-1));
        SIGNAL Multiplier85Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.577708,exponentBits,mantissaBits-1));
        SIGNAL Multiplier86Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.98124,exponentBits,mantissaBits-1));
        SIGNAL Multiplier88Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.960334,exponentBits,mantissaBits-1));
        SIGNAL Multiplier89Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.336149,exponentBits,mantissaBits-1));
        SIGNAL Multiplier90Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.99914,exponentBits,mantissaBits-1));
        SIGNAL Multiplier92Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.551341,exponentBits,mantissaBits-1));
        SIGNAL Multiplier93Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.926235,exponentBits,mantissaBits-1));
        SIGNAL Multiplier94Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.981519,exponentBits,mantissaBits-1));
        SIGNAL Multiplier95Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.989597,exponentBits,mantissaBits-1));
        SIGNAL Multiplier96Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.986786,exponentBits,mantissaBits-1));
        SIGNAL Multiplier97Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.995641,exponentBits,mantissaBits-1));
        SIGNAL Multiplier99Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.664315,exponentBits,mantissaBits-1));
        SIGNAL Multiplier101Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.634118,exponentBits,mantissaBits-1));
        SIGNAL Multiplier103Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.94312,exponentBits,mantissaBits-1));
        SIGNAL Multiplier105Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.970921,exponentBits,mantissaBits-1));
        SIGNAL Multiplier106Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.67214,exponentBits,mantissaBits-1));
        SIGNAL Multiplier108Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.98927,exponentBits,mantissaBits-1));
        SIGNAL Multiplier109Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.997554,exponentBits,mantissaBits-1));
        SIGNAL Multiplier110Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.414069,exponentBits,mantissaBits-1));
        SIGNAL Multiplier112Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.853307,exponentBits,mantissaBits-1));
        SIGNAL Multiplier113Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.886527,exponentBits,mantissaBits-1));
        SIGNAL Multiplier115Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.554692,exponentBits,mantissaBits-1));
        SIGNAL Multiplier116Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.989739,exponentBits,mantissaBits-1));
        SIGNAL Multiplier117Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.549861,exponentBits,mantissaBits-1));
        SIGNAL Multiplier120Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.994862,exponentBits,mantissaBits-1));
        SIGNAL Multiplier121Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.817897,exponentBits,mantissaBits-1));
        SIGNAL Multiplier122Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.912886,exponentBits,mantissaBits-1));
        SIGNAL Multiplier124Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.976301,exponentBits,mantissaBits-1));
        SIGNAL Multiplier125Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.98888,exponentBits,mantissaBits-1));
        SIGNAL Multiplier126Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.558577,exponentBits,mantissaBits-1));
        SIGNAL Multiplier128Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.731617,exponentBits,mantissaBits-1));
        SIGNAL Multiplier129Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.954043,exponentBits,mantissaBits-1));
        SIGNAL Multiplier131Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.646579,exponentBits,mantissaBits-1));
        SIGNAL Multiplier132Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.985013,exponentBits,mantissaBits-1));
        SIGNAL Multiplier133Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.592017,exponentBits,mantissaBits-1));
        SIGNAL Multiplier136Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.479802,exponentBits,mantissaBits-1));
        SIGNAL Multiplier138Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.927615,exponentBits,mantissaBits-1));
        SIGNAL Multiplier139Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.792795,exponentBits,mantissaBits-1));
        SIGNAL Multiplier141Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.907425,exponentBits,mantissaBits-1));
        SIGNAL Multiplier142Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.948402,exponentBits,mantissaBits-1));
        SIGNAL Multiplier143Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.83894,exponentBits,mantissaBits-1));
        SIGNAL Multiplier144Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.898142,exponentBits,mantissaBits-1));
        SIGNAL Multiplier146Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.826105,exponentBits,mantissaBits-1));
        SIGNAL Multiplier147Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.838083,exponentBits,mantissaBits-1));
        SIGNAL Multiplier149Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.970921,exponentBits,mantissaBits-1));
        SIGNAL Multiplier150Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.67214,exponentBits,mantissaBits-1));
        SIGNAL Multiplier152Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.98927,exponentBits,mantissaBits-1));
        SIGNAL Multiplier153Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.997554,exponentBits,mantissaBits-1));
        SIGNAL Multiplier154Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.414069,exponentBits,mantissaBits-1));
        SIGNAL Multiplier156Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.853307,exponentBits,mantissaBits-1));
        SIGNAL Multiplier157Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.886527,exponentBits,mantissaBits-1));
        SIGNAL Multiplier159Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.554692,exponentBits,mantissaBits-1));
        SIGNAL Multiplier160Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.989739,exponentBits,mantissaBits-1));
        SIGNAL Multiplier161Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.549861,exponentBits,mantissaBits-1));
        SIGNAL Multiplier164Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.970629,exponentBits,mantissaBits-1));
        SIGNAL Multiplier165Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.817897,exponentBits,mantissaBits-1));
        SIGNAL Multiplier166Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.912886,exponentBits,mantissaBits-1));
        SIGNAL Multiplier168Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.976301,exponentBits,mantissaBits-1));
        SIGNAL Multiplier169Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.98888,exponentBits,mantissaBits-1));
        SIGNAL Multiplier170Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.558577,exponentBits,mantissaBits-1));
        SIGNAL Multiplier172Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.731617,exponentBits,mantissaBits-1));
        SIGNAL Multiplier173Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.954043,exponentBits,mantissaBits-1));
        SIGNAL Multiplier175Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.646579,exponentBits,mantissaBits-1));
        SIGNAL Multiplier176Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.985013,exponentBits,mantissaBits-1));
        SIGNAL Multiplier177Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.592017,exponentBits,mantissaBits-1));
        SIGNAL Multiplier180Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.673404,exponentBits,mantissaBits-1));
        SIGNAL Multiplier182Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.750079,exponentBits,mantissaBits-1));
        SIGNAL Multiplier183Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.947231,exponentBits,mantissaBits-1));
        SIGNAL Multiplier185Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.907425,exponentBits,mantissaBits-1));
        SIGNAL Multiplier186Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.74707,exponentBits,mantissaBits-1));
        SIGNAL Multiplier187Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.617466,exponentBits,mantissaBits-1));
        SIGNAL Multiplier188Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.981367,exponentBits,mantissaBits-1));
        SIGNAL Multiplier190Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.826105,exponentBits,mantissaBits-1));
        SIGNAL Multiplier191Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.898792,exponentBits,mantissaBits-1));
        SIGNAL Multiplier194Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.995408,exponentBits,mantissaBits-1));
        SIGNAL Multiplier195Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.970921,exponentBits,mantissaBits-1));
        SIGNAL Multiplier196Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.67214,exponentBits,mantissaBits-1));
        SIGNAL Multiplier198Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.98927,exponentBits,mantissaBits-1));
        SIGNAL Multiplier199Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.966381,exponentBits,mantissaBits-1));
        SIGNAL Multiplier200Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.690672,exponentBits,mantissaBits-1));
        SIGNAL Multiplier202Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.853307,exponentBits,mantissaBits-1));
        SIGNAL Multiplier203Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.886527,exponentBits,mantissaBits-1));
        SIGNAL Multiplier205Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.554692,exponentBits,mantissaBits-1));
        SIGNAL Multiplier206Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.94187,exponentBits,mantissaBits-1));
        SIGNAL Multiplier207Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.763101,exponentBits,mantissaBits-1));
        SIGNAL Multiplier210Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.951966,exponentBits,mantissaBits-1));
        SIGNAL Multiplier211Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.817897,exponentBits,mantissaBits-1));
        SIGNAL Multiplier212Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.912886,exponentBits,mantissaBits-1));
        SIGNAL Multiplier214Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.976301,exponentBits,mantissaBits-1));
        SIGNAL Multiplier215Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.909585,exponentBits,mantissaBits-1));
        SIGNAL Multiplier216Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.82292,exponentBits,mantissaBits-1));
        SIGNAL Multiplier218Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.731617,exponentBits,mantissaBits-1));
        SIGNAL Multiplier219Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.954043,exponentBits,mantissaBits-1));
        SIGNAL Multiplier221Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.646579,exponentBits,mantissaBits-1));
        SIGNAL Multiplier222Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.790147,exponentBits,mantissaBits-1));
        SIGNAL Multiplier223Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.929014,exponentBits,mantissaBits-1));
        SIGNAL Multiplier226Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.7375,exponentBits,mantissaBits-1));
        SIGNAL Multiplier228Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.927615,exponentBits,mantissaBits-1));
        SIGNAL Multiplier229Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.792795,exponentBits,mantissaBits-1));
        SIGNAL Multiplier231Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.807766,exponentBits,mantissaBits-1));
        SIGNAL Multiplier232Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.907576,exponentBits,mantissaBits-1));
        SIGNAL Multiplier233Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.83894,exponentBits,mantissaBits-1));
        SIGNAL Multiplier234Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.898142,exponentBits,mantissaBits-1));
        SIGNAL Multiplier236Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.919167,exponentBits,mantissaBits-1));
        SIGNAL Multiplier237Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.781132,exponentBits,mantissaBits-1));
        SIGNAL Multiplier239Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.970921,exponentBits,mantissaBits-1));
        SIGNAL Multiplier240Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.67214,exponentBits,mantissaBits-1));
        SIGNAL Multiplier242Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.98927,exponentBits,mantissaBits-1));
        SIGNAL Multiplier243Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.966381,exponentBits,mantissaBits-1));
        SIGNAL Multiplier244Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.690672,exponentBits,mantissaBits-1));
        SIGNAL Multiplier246Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.853307,exponentBits,mantissaBits-1));
        SIGNAL Multiplier247Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.886527,exponentBits,mantissaBits-1));
        SIGNAL Multiplier249Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.554692,exponentBits,mantissaBits-1));
        SIGNAL Multiplier250Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.94187,exponentBits,mantissaBits-1));
        SIGNAL Multiplier251Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.763101,exponentBits,mantissaBits-1));
        SIGNAL Multiplier254Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.840616,exponentBits,mantissaBits-1));
        SIGNAL Multiplier255Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.817897,exponentBits,mantissaBits-1));
        SIGNAL Multiplier256Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.912886,exponentBits,mantissaBits-1));
        SIGNAL Multiplier258Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.976301,exponentBits,mantissaBits-1));
        SIGNAL Multiplier259Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.909585,exponentBits,mantissaBits-1));
        SIGNAL Multiplier260Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.82292,exponentBits,mantissaBits-1));
        SIGNAL Multiplier262Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.731617,exponentBits,mantissaBits-1));
        SIGNAL Multiplier263Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.954043,exponentBits,mantissaBits-1));
        SIGNAL Multiplier265Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.646579,exponentBits,mantissaBits-1));
        SIGNAL Multiplier266Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.790147,exponentBits,mantissaBits-1));
        SIGNAL Multiplier267Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.929014,exponentBits,mantissaBits-1));
        SIGNAL Multiplier270Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.896858,exponentBits,mantissaBits-1));
        SIGNAL Multiplier272Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.750079,exponentBits,mantissaBits-1));
        SIGNAL Multiplier273Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.947231,exponentBits,mantissaBits-1));
        SIGNAL Multiplier275Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.807766,exponentBits,mantissaBits-1));
        SIGNAL Multiplier276Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.825885,exponentBits,mantissaBits-1));
        SIGNAL Multiplier277Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.617466,exponentBits,mantissaBits-1));
        SIGNAL Multiplier278Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.981367,exponentBits,mantissaBits-1));
        SIGNAL Multiplier280Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.919167,exponentBits,mantissaBits-1));
        SIGNAL Multiplier281Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.93358,exponentBits,mantissaBits-1));
        SIGNAL Multiplier284Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.469245,exponentBits,mantissaBits-1));
        SIGNAL Multiplier286Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.848299,exponentBits,mantissaBits-1));
        SIGNAL Multiplier287Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.895308,exponentBits,mantissaBits-1));
        SIGNAL Multiplier288Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.842608,exponentBits,mantissaBits-1));
        SIGNAL Multiplier290Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870697,exponentBits,mantissaBits-1));
        SIGNAL Multiplier291Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.945793,exponentBits,mantissaBits-1));
        SIGNAL Multiplier292Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.95487,exponentBits,mantissaBits-1));
        SIGNAL Multiplier293Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870404,exponentBits,mantissaBits-1));
        SIGNAL Multiplier294Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.780732,exponentBits,mantissaBits-1));
        SIGNAL Multiplier295Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.810846,exponentBits,mantissaBits-1));
        SIGNAL Multiplier297Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.991361,exponentBits,mantissaBits-1));
        SIGNAL Multiplier298Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.669241,exponentBits,mantissaBits-1));
        SIGNAL Multiplier299Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.97158,exponentBits,mantissaBits-1));
        SIGNAL Multiplier301Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870697,exponentBits,mantissaBits-1));
        SIGNAL Multiplier302Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.75369,exponentBits,mantissaBits-1));
        SIGNAL Multiplier303Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.77448,exponentBits,mantissaBits-1));
        SIGNAL Multiplier304Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870404,exponentBits,mantissaBits-1));
        SIGNAL Multiplier305Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.933776,exponentBits,mantissaBits-1));
        SIGNAL Multiplier306Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.660973,exponentBits,mantissaBits-1));
        SIGNAL Multiplier308Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870239,exponentBits,mantissaBits-1));
        SIGNAL Multiplier310Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.756327,exponentBits,mantissaBits-1));
        SIGNAL Multiplier311Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.890735,exponentBits,mantissaBits-1));
        SIGNAL Multiplier312Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.689002,exponentBits,mantissaBits-1));
        SIGNAL Multiplier313Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.966814,exponentBits,mantissaBits-1));
        SIGNAL Multiplier315Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.551341,exponentBits,mantissaBits-1));
        SIGNAL Multiplier316Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.795357,exponentBits,mantissaBits-1));
        SIGNAL Multiplier317Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.746308,exponentBits,mantissaBits-1));
        SIGNAL Multiplier318Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.989597,exponentBits,mantissaBits-1));
        SIGNAL Multiplier319Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.577708,exponentBits,mantissaBits-1));
        SIGNAL Multiplier320Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.618274,exponentBits,mantissaBits-1));
        SIGNAL Multiplier322Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.952809,exponentBits,mantissaBits-1));
        SIGNAL Multiplier323Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.495915,exponentBits,mantissaBits-1));
        SIGNAL Multiplier324Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.993928,exponentBits,mantissaBits-1));
        SIGNAL Multiplier326Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.551341,exponentBits,mantissaBits-1));
        SIGNAL Multiplier327Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.926235,exponentBits,mantissaBits-1));
        SIGNAL Multiplier328Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.616494,exponentBits,mantissaBits-1));
        SIGNAL Multiplier329Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.989597,exponentBits,mantissaBits-1));
        SIGNAL Multiplier330Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.986786,exponentBits,mantissaBits-1));
        SIGNAL Multiplier331Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.464416,exponentBits,mantissaBits-1));
        SIGNAL Multiplier333Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.770987,exponentBits,mantissaBits-1));
        SIGNAL Multiplier335Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.906302,exponentBits,mantissaBits-1));
        SIGNAL Multiplier337Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.800117,exponentBits,mantissaBits-1));
        SIGNAL Multiplier338Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.848299,exponentBits,mantissaBits-1));
        SIGNAL Multiplier339Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.562709,exponentBits,mantissaBits-1));
        SIGNAL Multiplier340Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.988453,exponentBits,mantissaBits-1));
        SIGNAL Multiplier342Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870697,exponentBits,mantissaBits-1));
        SIGNAL Multiplier343Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.945793,exponentBits,mantissaBits-1));
        SIGNAL Multiplier344Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.729204,exponentBits,mantissaBits-1));
        SIGNAL Multiplier345Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870404,exponentBits,mantissaBits-1));
        SIGNAL Multiplier346Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.780732,exponentBits,mantissaBits-1));
        SIGNAL Multiplier347Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.917308,exponentBits,mantissaBits-1));
        SIGNAL Multiplier349Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.979033,exponentBits,mantissaBits-1));
        SIGNAL Multiplier350Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.453222,exponentBits,mantissaBits-1));
        SIGNAL Multiplier351Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.996146,exponentBits,mantissaBits-1));
        SIGNAL Multiplier353Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870697,exponentBits,mantissaBits-1));
        SIGNAL Multiplier354Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.75369,exponentBits,mantissaBits-1));
        SIGNAL Multiplier355Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.936763,exponentBits,mantissaBits-1));
        SIGNAL Multiplier356Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870404,exponentBits,mantissaBits-1));
        SIGNAL Multiplier357Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.933776,exponentBits,mantissaBits-1));
        SIGNAL Multiplier358Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.973389,exponentBits,mantissaBits-1));
        SIGNAL Multiplier360Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.818419,exponentBits,mantissaBits-1));
        SIGNAL Multiplier362Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.940496,exponentBits,mantissaBits-1));
        SIGNAL Multiplier363Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.890735,exponentBits,mantissaBits-1));
        SIGNAL Multiplier364Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.382644,exponentBits,mantissaBits-1));
        SIGNAL Multiplier365Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.998354,exponentBits,mantissaBits-1));
        SIGNAL Multiplier367Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.551341,exponentBits,mantissaBits-1));
        SIGNAL Multiplier368Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.795357,exponentBits,mantissaBits-1));
        SIGNAL Multiplier369Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.948695,exponentBits,mantissaBits-1));
        SIGNAL Multiplier370Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.989597,exponentBits,mantissaBits-1));
        SIGNAL Multiplier371Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.577708,exponentBits,mantissaBits-1));
        SIGNAL Multiplier372Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.98124,exponentBits,mantissaBits-1));
        SIGNAL Multiplier374Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.960334,exponentBits,mantissaBits-1));
        SIGNAL Multiplier375Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.336149,exponentBits,mantissaBits-1));
        SIGNAL Multiplier376Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.99914,exponentBits,mantissaBits-1));
        SIGNAL Multiplier378Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.551341,exponentBits,mantissaBits-1));
        SIGNAL Multiplier379Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.926235,exponentBits,mantissaBits-1));
        SIGNAL Multiplier380Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.981519,exponentBits,mantissaBits-1));
        SIGNAL Multiplier381Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.989597,exponentBits,mantissaBits-1));
        SIGNAL Multiplier382Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.986786,exponentBits,mantissaBits-1));
        SIGNAL Multiplier383Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.995641,exponentBits,mantissaBits-1));
        SIGNAL Multiplier385Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.664315,exponentBits,mantissaBits-1));
        SIGNAL Multiplier387Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.978597,exponentBits,mantissaBits-1));
        SIGNAL Multiplier389Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.655866,exponentBits,mantissaBits-1));
        SIGNAL Multiplier391Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.970921,exponentBits,mantissaBits-1));
        SIGNAL Multiplier392Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.67214,exponentBits,mantissaBits-1));
        SIGNAL Multiplier394Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.98927,exponentBits,mantissaBits-1));
        SIGNAL Multiplier395Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.997554,exponentBits,mantissaBits-1));
        SIGNAL Multiplier396Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.414069,exponentBits,mantissaBits-1));
        SIGNAL Multiplier398Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.853307,exponentBits,mantissaBits-1));
        SIGNAL Multiplier399Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.886527,exponentBits,mantissaBits-1));
        SIGNAL Multiplier401Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.554692,exponentBits,mantissaBits-1));
        SIGNAL Multiplier402Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.989739,exponentBits,mantissaBits-1));
        SIGNAL Multiplier403Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.549861,exponentBits,mantissaBits-1));
        SIGNAL Multiplier406Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.994862,exponentBits,mantissaBits-1));
        SIGNAL Multiplier407Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.817897,exponentBits,mantissaBits-1));
        SIGNAL Multiplier408Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.912886,exponentBits,mantissaBits-1));
        SIGNAL Multiplier410Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.976301,exponentBits,mantissaBits-1));
        SIGNAL Multiplier411Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.98888,exponentBits,mantissaBits-1));
        SIGNAL Multiplier412Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.558577,exponentBits,mantissaBits-1));
        SIGNAL Multiplier414Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.731617,exponentBits,mantissaBits-1));
        SIGNAL Multiplier415Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.954043,exponentBits,mantissaBits-1));
        SIGNAL Multiplier417Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.646579,exponentBits,mantissaBits-1));
        SIGNAL Multiplier418Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.985013,exponentBits,mantissaBits-1));
        SIGNAL Multiplier419Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.592017,exponentBits,mantissaBits-1));
        SIGNAL Multiplier422Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.479802,exponentBits,mantissaBits-1));
        SIGNAL Multiplier424Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.927615,exponentBits,mantissaBits-1));
        SIGNAL Multiplier425Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.792795,exponentBits,mantissaBits-1));
        SIGNAL Multiplier427Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.907425,exponentBits,mantissaBits-1));
        SIGNAL Multiplier428Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.948402,exponentBits,mantissaBits-1));
        SIGNAL Multiplier429Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.83894,exponentBits,mantissaBits-1));
        SIGNAL Multiplier430Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.898142,exponentBits,mantissaBits-1));
        SIGNAL Multiplier432Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.826105,exponentBits,mantissaBits-1));
        SIGNAL Multiplier433Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.838083,exponentBits,mantissaBits-1));
        SIGNAL Multiplier435Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.970921,exponentBits,mantissaBits-1));
        SIGNAL Multiplier436Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.67214,exponentBits,mantissaBits-1));
        SIGNAL Multiplier438Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.98927,exponentBits,mantissaBits-1));
        SIGNAL Multiplier439Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.997554,exponentBits,mantissaBits-1));
        SIGNAL Multiplier440Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.414069,exponentBits,mantissaBits-1));
        SIGNAL Multiplier442Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.853307,exponentBits,mantissaBits-1));
        SIGNAL Multiplier443Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.886527,exponentBits,mantissaBits-1));
        SIGNAL Multiplier445Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.554692,exponentBits,mantissaBits-1));
        SIGNAL Multiplier446Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.989739,exponentBits,mantissaBits-1));
        SIGNAL Multiplier447Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.549861,exponentBits,mantissaBits-1));
        SIGNAL Multiplier450Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.970629,exponentBits,mantissaBits-1));
        SIGNAL Multiplier451Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.817897,exponentBits,mantissaBits-1));
        SIGNAL Multiplier452Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.912886,exponentBits,mantissaBits-1));
        SIGNAL Multiplier454Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.976301,exponentBits,mantissaBits-1));
        SIGNAL Multiplier455Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.98888,exponentBits,mantissaBits-1));
        SIGNAL Multiplier456Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.558577,exponentBits,mantissaBits-1));
        SIGNAL Multiplier458Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.731617,exponentBits,mantissaBits-1));
        SIGNAL Multiplier459Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.954043,exponentBits,mantissaBits-1));
        SIGNAL Multiplier461Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.646579,exponentBits,mantissaBits-1));
        SIGNAL Multiplier462Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.985013,exponentBits,mantissaBits-1));
        SIGNAL Multiplier463Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.592017,exponentBits,mantissaBits-1));
        SIGNAL Multiplier466Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.673404,exponentBits,mantissaBits-1));
        SIGNAL Multiplier468Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.750079,exponentBits,mantissaBits-1));
        SIGNAL Multiplier469Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.947231,exponentBits,mantissaBits-1));
        SIGNAL Multiplier471Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.907425,exponentBits,mantissaBits-1));
        SIGNAL Multiplier472Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.74707,exponentBits,mantissaBits-1));
        SIGNAL Multiplier473Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.617466,exponentBits,mantissaBits-1));
        SIGNAL Multiplier474Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.981367,exponentBits,mantissaBits-1));
        SIGNAL Multiplier476Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.826105,exponentBits,mantissaBits-1));
        SIGNAL Multiplier477Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.898792,exponentBits,mantissaBits-1));
        SIGNAL Multiplier480Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.935776,exponentBits,mantissaBits-1));
        SIGNAL Multiplier481Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.970921,exponentBits,mantissaBits-1));
        SIGNAL Multiplier482Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.67214,exponentBits,mantissaBits-1));
        SIGNAL Multiplier484Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.98927,exponentBits,mantissaBits-1));
        SIGNAL Multiplier485Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.966381,exponentBits,mantissaBits-1));
        SIGNAL Multiplier486Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.690672,exponentBits,mantissaBits-1));
        SIGNAL Multiplier488Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.853307,exponentBits,mantissaBits-1));
        SIGNAL Multiplier489Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.886527,exponentBits,mantissaBits-1));
        SIGNAL Multiplier491Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.554692,exponentBits,mantissaBits-1));
        SIGNAL Multiplier492Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.94187,exponentBits,mantissaBits-1));
        SIGNAL Multiplier493Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.763101,exponentBits,mantissaBits-1));
        SIGNAL Multiplier496Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.951966,exponentBits,mantissaBits-1));
        SIGNAL Multiplier497Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.817897,exponentBits,mantissaBits-1));
        SIGNAL Multiplier498Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.912886,exponentBits,mantissaBits-1));
        SIGNAL Multiplier500Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.976301,exponentBits,mantissaBits-1));
        SIGNAL Multiplier501Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.909585,exponentBits,mantissaBits-1));
        SIGNAL Multiplier502Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.82292,exponentBits,mantissaBits-1));
        SIGNAL Multiplier504Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.731617,exponentBits,mantissaBits-1));
        SIGNAL Multiplier505Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.954043,exponentBits,mantissaBits-1));
        SIGNAL Multiplier507Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.646579,exponentBits,mantissaBits-1));
        SIGNAL Multiplier508Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.790147,exponentBits,mantissaBits-1));
        SIGNAL Multiplier509Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.929014,exponentBits,mantissaBits-1));
        SIGNAL Multiplier512Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.7375,exponentBits,mantissaBits-1));
        SIGNAL Multiplier514Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.927615,exponentBits,mantissaBits-1));
        SIGNAL Multiplier515Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.792795,exponentBits,mantissaBits-1));
        SIGNAL Multiplier517Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.807766,exponentBits,mantissaBits-1));
        SIGNAL Multiplier518Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.907576,exponentBits,mantissaBits-1));
        SIGNAL Multiplier519Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.83894,exponentBits,mantissaBits-1));
        SIGNAL Multiplier520Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.898142,exponentBits,mantissaBits-1));
        SIGNAL Multiplier522Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.919167,exponentBits,mantissaBits-1));
        SIGNAL Multiplier523Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.781132,exponentBits,mantissaBits-1));
        SIGNAL Multiplier525Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.970921,exponentBits,mantissaBits-1));
        SIGNAL Multiplier526Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.67214,exponentBits,mantissaBits-1));
        SIGNAL Multiplier528Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.98927,exponentBits,mantissaBits-1));
        SIGNAL Multiplier529Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.966381,exponentBits,mantissaBits-1));
        SIGNAL Multiplier530Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.690672,exponentBits,mantissaBits-1));
        SIGNAL Multiplier532Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.853307,exponentBits,mantissaBits-1));
        SIGNAL Multiplier533Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.886527,exponentBits,mantissaBits-1));
        SIGNAL Multiplier535Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.554692,exponentBits,mantissaBits-1));
        SIGNAL Multiplier536Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.94187,exponentBits,mantissaBits-1));
        SIGNAL Multiplier537Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.763101,exponentBits,mantissaBits-1));
        SIGNAL Multiplier540Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.840616,exponentBits,mantissaBits-1));
        SIGNAL Multiplier541Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.817897,exponentBits,mantissaBits-1));
        SIGNAL Multiplier542Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.912886,exponentBits,mantissaBits-1));
        SIGNAL Multiplier544Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.976301,exponentBits,mantissaBits-1));
        SIGNAL Multiplier545Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.909585,exponentBits,mantissaBits-1));
        SIGNAL Multiplier546Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.82292,exponentBits,mantissaBits-1));
        SIGNAL Multiplier548Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.731617,exponentBits,mantissaBits-1));
        SIGNAL Multiplier549Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.954043,exponentBits,mantissaBits-1));
        SIGNAL Multiplier551Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.646579,exponentBits,mantissaBits-1));
        SIGNAL Multiplier552Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.790147,exponentBits,mantissaBits-1));
        SIGNAL Multiplier553Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.929014,exponentBits,mantissaBits-1));
        SIGNAL Multiplier556Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.896858,exponentBits,mantissaBits-1));
        SIGNAL Multiplier558Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.750079,exponentBits,mantissaBits-1));
        SIGNAL Multiplier559Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.947231,exponentBits,mantissaBits-1));
        SIGNAL Multiplier561Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.807766,exponentBits,mantissaBits-1));
        SIGNAL Multiplier562Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.825885,exponentBits,mantissaBits-1));
        SIGNAL Multiplier563Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.617466,exponentBits,mantissaBits-1));
        SIGNAL Multiplier564Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.981367,exponentBits,mantissaBits-1));
        SIGNAL Multiplier566Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.919167,exponentBits,mantissaBits-1));
        SIGNAL Multiplier567Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.93358,exponentBits,mantissaBits-1));
        SIGNAL Multiplier570Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.776577,exponentBits,mantissaBits-1));
        SIGNAL Multiplier573Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.848299,exponentBits,mantissaBits-1));
        SIGNAL Multiplier574Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.895308,exponentBits,mantissaBits-1));
        SIGNAL Multiplier575Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.842608,exponentBits,mantissaBits-1));
        SIGNAL Multiplier577Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870697,exponentBits,mantissaBits-1));
        SIGNAL Multiplier578Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.945793,exponentBits,mantissaBits-1));
        SIGNAL Multiplier579Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.95487,exponentBits,mantissaBits-1));
        SIGNAL Multiplier580Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870404,exponentBits,mantissaBits-1));
        SIGNAL Multiplier581Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.780732,exponentBits,mantissaBits-1));
        SIGNAL Multiplier582Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.810846,exponentBits,mantissaBits-1));
        SIGNAL Multiplier584Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.531606,exponentBits,mantissaBits-1));
        SIGNAL Multiplier585Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.669241,exponentBits,mantissaBits-1));
        SIGNAL Multiplier586Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.97158,exponentBits,mantissaBits-1));
        SIGNAL Multiplier588Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870697,exponentBits,mantissaBits-1));
        SIGNAL Multiplier589Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.75369,exponentBits,mantissaBits-1));
        SIGNAL Multiplier590Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.77448,exponentBits,mantissaBits-1));
        SIGNAL Multiplier591Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870404,exponentBits,mantissaBits-1));
        SIGNAL Multiplier592Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.933776,exponentBits,mantissaBits-1));
        SIGNAL Multiplier593Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.660973,exponentBits,mantissaBits-1));
        SIGNAL Multiplier595Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870862,exponentBits,mantissaBits-1));
        SIGNAL Multiplier597Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.85073,exponentBits,mantissaBits-1));
        SIGNAL Multiplier598Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.890735,exponentBits,mantissaBits-1));
        SIGNAL Multiplier599Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.689002,exponentBits,mantissaBits-1));
        SIGNAL Multiplier600Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.966814,exponentBits,mantissaBits-1));
        SIGNAL Multiplier602Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.551341,exponentBits,mantissaBits-1));
        SIGNAL Multiplier603Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.795357,exponentBits,mantissaBits-1));
        SIGNAL Multiplier604Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.746308,exponentBits,mantissaBits-1));
        SIGNAL Multiplier605Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.989597,exponentBits,mantissaBits-1));
        SIGNAL Multiplier606Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.577708,exponentBits,mantissaBits-1));
        SIGNAL Multiplier607Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.618274,exponentBits,mantissaBits-1));
        SIGNAL Multiplier609Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.735141,exponentBits,mantissaBits-1));
        SIGNAL Multiplier610Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.495915,exponentBits,mantissaBits-1));
        SIGNAL Multiplier611Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.993928,exponentBits,mantissaBits-1));
        SIGNAL Multiplier613Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.551341,exponentBits,mantissaBits-1));
        SIGNAL Multiplier614Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.926235,exponentBits,mantissaBits-1));
        SIGNAL Multiplier615Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.616494,exponentBits,mantissaBits-1));
        SIGNAL Multiplier616Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.989597,exponentBits,mantissaBits-1));
        SIGNAL Multiplier617Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.986786,exponentBits,mantissaBits-1));
        SIGNAL Multiplier618Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.464416,exponentBits,mantissaBits-1));
        SIGNAL Multiplier620Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.938375,exponentBits,mantissaBits-1));
        SIGNAL Multiplier622Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.635106,exponentBits,mantissaBits-1));
        SIGNAL Multiplier624Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.969587,exponentBits,mantissaBits-1));
        SIGNAL Multiplier625Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.848299,exponentBits,mantissaBits-1));
        SIGNAL Multiplier626Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.562709,exponentBits,mantissaBits-1));
        SIGNAL Multiplier627Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.988453,exponentBits,mantissaBits-1));
        SIGNAL Multiplier629Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870697,exponentBits,mantissaBits-1));
        SIGNAL Multiplier630Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.945793,exponentBits,mantissaBits-1));
        SIGNAL Multiplier631Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.729204,exponentBits,mantissaBits-1));
        SIGNAL Multiplier632Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870404,exponentBits,mantissaBits-1));
        SIGNAL Multiplier633Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.780732,exponentBits,mantissaBits-1));
        SIGNAL Multiplier634Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.917308,exponentBits,mantissaBits-1));
        SIGNAL Multiplier636Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.631626,exponentBits,mantissaBits-1));
        SIGNAL Multiplier637Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.453222,exponentBits,mantissaBits-1));
        SIGNAL Multiplier638Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.996146,exponentBits,mantissaBits-1));
        SIGNAL Multiplier640Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870697,exponentBits,mantissaBits-1));
        SIGNAL Multiplier641Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.75369,exponentBits,mantissaBits-1));
        SIGNAL Multiplier642Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.936763,exponentBits,mantissaBits-1));
        SIGNAL Multiplier643Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870404,exponentBits,mantissaBits-1));
        SIGNAL Multiplier644Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.933776,exponentBits,mantissaBits-1));
        SIGNAL Multiplier645Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.973389,exponentBits,mantissaBits-1));
        SIGNAL Multiplier647Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.912549,exponentBits,mantissaBits-1));
        SIGNAL Multiplier649Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.658116,exponentBits,mantissaBits-1));
        SIGNAL Multiplier650Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.890735,exponentBits,mantissaBits-1));
        SIGNAL Multiplier651Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.382644,exponentBits,mantissaBits-1));
        SIGNAL Multiplier652Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.998354,exponentBits,mantissaBits-1));
        SIGNAL Multiplier654Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.551341,exponentBits,mantissaBits-1));
        SIGNAL Multiplier655Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.795357,exponentBits,mantissaBits-1));
        SIGNAL Multiplier656Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.948695,exponentBits,mantissaBits-1));
        SIGNAL Multiplier657Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.989597,exponentBits,mantissaBits-1));
        SIGNAL Multiplier658Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.577708,exponentBits,mantissaBits-1));
        SIGNAL Multiplier659Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.98124,exponentBits,mantissaBits-1));
        SIGNAL Multiplier661Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.712179,exponentBits,mantissaBits-1));
        SIGNAL Multiplier662Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.336149,exponentBits,mantissaBits-1));
        SIGNAL Multiplier663Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.99914,exponentBits,mantissaBits-1));
        SIGNAL Multiplier665Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.551341,exponentBits,mantissaBits-1));
        SIGNAL Multiplier666Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.926235,exponentBits,mantissaBits-1));
        SIGNAL Multiplier667Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.981519,exponentBits,mantissaBits-1));
        SIGNAL Multiplier668Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.989597,exponentBits,mantissaBits-1));
        SIGNAL Multiplier669Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.986786,exponentBits,mantissaBits-1));
        SIGNAL Multiplier670Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.995641,exponentBits,mantissaBits-1));
        SIGNAL Multiplier672Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.97267,exponentBits,mantissaBits-1));
        SIGNAL Multiplier674Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.53135,exponentBits,mantissaBits-1));
        SIGNAL Multiplier676Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.913608,exponentBits,mantissaBits-1));
        SIGNAL Multiplier678Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.965849,exponentBits,mantissaBits-1));
        SIGNAL Multiplier679Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.692695,exponentBits,mantissaBits-1));
        SIGNAL Multiplier681Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.880399,exponentBits,mantissaBits-1));
        SIGNAL Multiplier682Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.997554,exponentBits,mantissaBits-1));
        SIGNAL Multiplier683Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.414069,exponentBits,mantissaBits-1));
        SIGNAL Multiplier685Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.91966,exponentBits,mantissaBits-1));
        SIGNAL Multiplier686Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.806938,exponentBits,mantissaBits-1));
        SIGNAL Multiplier688Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.860235,exponentBits,mantissaBits-1));
        SIGNAL Multiplier689Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.989739,exponentBits,mantissaBits-1));
        SIGNAL Multiplier690Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.549861,exponentBits,mantissaBits-1));
        SIGNAL Multiplier693Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.984104,exponentBits,mantissaBits-1));
        SIGNAL Multiplier694Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.793165,exponentBits,mantissaBits-1));
        SIGNAL Multiplier695Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.927417,exponentBits,mantissaBits-1));
        SIGNAL Multiplier697Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.726095,exponentBits,mantissaBits-1));
        SIGNAL Multiplier698Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.98888,exponentBits,mantissaBits-1));
        SIGNAL Multiplier699Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.558577,exponentBits,mantissaBits-1));
        SIGNAL Multiplier701Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.649155,exponentBits,mantissaBits-1));
        SIGNAL Multiplier702Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.975801,exponentBits,mantissaBits-1));
        SIGNAL Multiplier704Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.955917,exponentBits,mantissaBits-1));
        SIGNAL Multiplier705Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.985013,exponentBits,mantissaBits-1));
        SIGNAL Multiplier706Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.592017,exponentBits,mantissaBits-1));
        SIGNAL Multiplier709Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.598812,exponentBits,mantissaBits-1));
        SIGNAL Multiplier711Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.927615,exponentBits,mantissaBits-1));
        SIGNAL Multiplier712Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.792795,exponentBits,mantissaBits-1));
        SIGNAL Multiplier714Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.907425,exponentBits,mantissaBits-1));
        SIGNAL Multiplier715Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.948402,exponentBits,mantissaBits-1));
        SIGNAL Multiplier716Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.83894,exponentBits,mantissaBits-1));
        SIGNAL Multiplier717Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.898142,exponentBits,mantissaBits-1));
        SIGNAL Multiplier719Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.826105,exponentBits,mantissaBits-1));
        SIGNAL Multiplier720Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.838083,exponentBits,mantissaBits-1));
        SIGNAL Multiplier722Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.965849,exponentBits,mantissaBits-1));
        SIGNAL Multiplier723Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.692695,exponentBits,mantissaBits-1));
        SIGNAL Multiplier725Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.880399,exponentBits,mantissaBits-1));
        SIGNAL Multiplier726Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.997554,exponentBits,mantissaBits-1));
        SIGNAL Multiplier727Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.414069,exponentBits,mantissaBits-1));
        SIGNAL Multiplier729Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.91966,exponentBits,mantissaBits-1));
        SIGNAL Multiplier730Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.806938,exponentBits,mantissaBits-1));
        SIGNAL Multiplier732Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.860235,exponentBits,mantissaBits-1));
        SIGNAL Multiplier733Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.989739,exponentBits,mantissaBits-1));
        SIGNAL Multiplier734Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.549861,exponentBits,mantissaBits-1));
        SIGNAL Multiplier737Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.932937,exponentBits,mantissaBits-1));
        SIGNAL Multiplier738Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.793165,exponentBits,mantissaBits-1));
        SIGNAL Multiplier739Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.927417,exponentBits,mantissaBits-1));
        SIGNAL Multiplier741Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.726095,exponentBits,mantissaBits-1));
        SIGNAL Multiplier742Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.98888,exponentBits,mantissaBits-1));
        SIGNAL Multiplier743Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.558577,exponentBits,mantissaBits-1));
        SIGNAL Multiplier745Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.649155,exponentBits,mantissaBits-1));
        SIGNAL Multiplier746Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.975801,exponentBits,mantissaBits-1));
        SIGNAL Multiplier748Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.955917,exponentBits,mantissaBits-1));
        SIGNAL Multiplier749Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.985013,exponentBits,mantissaBits-1));
        SIGNAL Multiplier750Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.592017,exponentBits,mantissaBits-1));
        SIGNAL Multiplier753Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.782438,exponentBits,mantissaBits-1));
        SIGNAL Multiplier755Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.750079,exponentBits,mantissaBits-1));
        SIGNAL Multiplier756Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.947231,exponentBits,mantissaBits-1));
        SIGNAL Multiplier758Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.907425,exponentBits,mantissaBits-1));
        SIGNAL Multiplier759Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.74707,exponentBits,mantissaBits-1));
        SIGNAL Multiplier760Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.617466,exponentBits,mantissaBits-1));
        SIGNAL Multiplier761Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.981367,exponentBits,mantissaBits-1));
        SIGNAL Multiplier763Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.826105,exponentBits,mantissaBits-1));
        SIGNAL Multiplier764Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.898792,exponentBits,mantissaBits-1));
        SIGNAL Multiplier767Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.987852,exponentBits,mantissaBits-1));
        SIGNAL Multiplier768Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.965849,exponentBits,mantissaBits-1));
        SIGNAL Multiplier769Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.692695,exponentBits,mantissaBits-1));
        SIGNAL Multiplier771Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.880399,exponentBits,mantissaBits-1));
        SIGNAL Multiplier772Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.966381,exponentBits,mantissaBits-1));
        SIGNAL Multiplier773Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.690672,exponentBits,mantissaBits-1));
        SIGNAL Multiplier775Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.91966,exponentBits,mantissaBits-1));
        SIGNAL Multiplier776Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.806938,exponentBits,mantissaBits-1));
        SIGNAL Multiplier778Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.860235,exponentBits,mantissaBits-1));
        SIGNAL Multiplier779Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.94187,exponentBits,mantissaBits-1));
        SIGNAL Multiplier780Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.763101,exponentBits,mantissaBits-1));
        SIGNAL Multiplier783Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.924413,exponentBits,mantissaBits-1));
        SIGNAL Multiplier784Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.793165,exponentBits,mantissaBits-1));
        SIGNAL Multiplier785Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.927417,exponentBits,mantissaBits-1));
        SIGNAL Multiplier787Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.726095,exponentBits,mantissaBits-1));
        SIGNAL Multiplier788Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.909585,exponentBits,mantissaBits-1));
        SIGNAL Multiplier789Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.82292,exponentBits,mantissaBits-1));
        SIGNAL Multiplier791Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.649155,exponentBits,mantissaBits-1));
        SIGNAL Multiplier792Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.975801,exponentBits,mantissaBits-1));
        SIGNAL Multiplier794Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.955917,exponentBits,mantissaBits-1));
        SIGNAL Multiplier795Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.790147,exponentBits,mantissaBits-1));
        SIGNAL Multiplier796Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.929014,exponentBits,mantissaBits-1));
        SIGNAL Multiplier799Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.798666,exponentBits,mantissaBits-1));
        SIGNAL Multiplier801Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.927615,exponentBits,mantissaBits-1));
        SIGNAL Multiplier802Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.792795,exponentBits,mantissaBits-1));
        SIGNAL Multiplier804Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.807766,exponentBits,mantissaBits-1));
        SIGNAL Multiplier805Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.907576,exponentBits,mantissaBits-1));
        SIGNAL Multiplier806Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.83894,exponentBits,mantissaBits-1));
        SIGNAL Multiplier807Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.898142,exponentBits,mantissaBits-1));
        SIGNAL Multiplier809Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.919167,exponentBits,mantissaBits-1));
        SIGNAL Multiplier810Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.781132,exponentBits,mantissaBits-1));
        SIGNAL Multiplier812Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.965849,exponentBits,mantissaBits-1));
        SIGNAL Multiplier813Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.692695,exponentBits,mantissaBits-1));
        SIGNAL Multiplier815Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.880399,exponentBits,mantissaBits-1));
        SIGNAL Multiplier816Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.966381,exponentBits,mantissaBits-1));
        SIGNAL Multiplier817Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.690672,exponentBits,mantissaBits-1));
        SIGNAL Multiplier819Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.91966,exponentBits,mantissaBits-1));
        SIGNAL Multiplier820Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.806938,exponentBits,mantissaBits-1));
        SIGNAL Multiplier822Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.860235,exponentBits,mantissaBits-1));
        SIGNAL Multiplier823Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.94187,exponentBits,mantissaBits-1));
        SIGNAL Multiplier824Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.763101,exponentBits,mantissaBits-1));
        SIGNAL Multiplier827Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.693688,exponentBits,mantissaBits-1));
        SIGNAL Multiplier828Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.793165,exponentBits,mantissaBits-1));
        SIGNAL Multiplier829Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.927417,exponentBits,mantissaBits-1));
        SIGNAL Multiplier831Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.726095,exponentBits,mantissaBits-1));
        SIGNAL Multiplier832Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.909585,exponentBits,mantissaBits-1));
        SIGNAL Multiplier833Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.82292,exponentBits,mantissaBits-1));
        SIGNAL Multiplier835Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.649155,exponentBits,mantissaBits-1));
        SIGNAL Multiplier836Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.975801,exponentBits,mantissaBits-1));
        SIGNAL Multiplier838Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.955917,exponentBits,mantissaBits-1));
        SIGNAL Multiplier839Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.790147,exponentBits,mantissaBits-1));
        SIGNAL Multiplier840Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.929014,exponentBits,mantissaBits-1));
        SIGNAL Multiplier843Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.965586,exponentBits,mantissaBits-1));
        SIGNAL Multiplier845Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.750079,exponentBits,mantissaBits-1));
        SIGNAL Multiplier846Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.947231,exponentBits,mantissaBits-1));
        SIGNAL Multiplier848Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.807766,exponentBits,mantissaBits-1));
        SIGNAL Multiplier849Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.825885,exponentBits,mantissaBits-1));
        SIGNAL Multiplier850Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.617466,exponentBits,mantissaBits-1));
        SIGNAL Multiplier851Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.981367,exponentBits,mantissaBits-1));
        SIGNAL Multiplier853Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.919167,exponentBits,mantissaBits-1));
        SIGNAL Multiplier854Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.93358,exponentBits,mantissaBits-1));
        SIGNAL Multiplier857Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.568305,exponentBits,mantissaBits-1));
        SIGNAL Multiplier859Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.848299,exponentBits,mantissaBits-1));
        SIGNAL Multiplier860Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.895308,exponentBits,mantissaBits-1));
        SIGNAL Multiplier861Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.842608,exponentBits,mantissaBits-1));
        SIGNAL Multiplier863Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870697,exponentBits,mantissaBits-1));
        SIGNAL Multiplier864Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.945793,exponentBits,mantissaBits-1));
        SIGNAL Multiplier865Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.95487,exponentBits,mantissaBits-1));
        SIGNAL Multiplier866Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870404,exponentBits,mantissaBits-1));
        SIGNAL Multiplier867Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.780732,exponentBits,mantissaBits-1));
        SIGNAL Multiplier868Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.810846,exponentBits,mantissaBits-1));
        SIGNAL Multiplier870Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.531606,exponentBits,mantissaBits-1));
        SIGNAL Multiplier871Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.669241,exponentBits,mantissaBits-1));
        SIGNAL Multiplier872Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.97158,exponentBits,mantissaBits-1));
        SIGNAL Multiplier874Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870697,exponentBits,mantissaBits-1));
        SIGNAL Multiplier875Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.75369,exponentBits,mantissaBits-1));
        SIGNAL Multiplier876Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.77448,exponentBits,mantissaBits-1));
        SIGNAL Multiplier877Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870404,exponentBits,mantissaBits-1));
        SIGNAL Multiplier878Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.933776,exponentBits,mantissaBits-1));
        SIGNAL Multiplier879Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.660973,exponentBits,mantissaBits-1));
        SIGNAL Multiplier881Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870862,exponentBits,mantissaBits-1));
        SIGNAL Multiplier883Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.888715,exponentBits,mantissaBits-1));
        SIGNAL Multiplier884Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.890735,exponentBits,mantissaBits-1));
        SIGNAL Multiplier885Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.689002,exponentBits,mantissaBits-1));
        SIGNAL Multiplier886Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.966814,exponentBits,mantissaBits-1));
        SIGNAL Multiplier888Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.551341,exponentBits,mantissaBits-1));
        SIGNAL Multiplier889Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.795357,exponentBits,mantissaBits-1));
        SIGNAL Multiplier890Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.746308,exponentBits,mantissaBits-1));
        SIGNAL Multiplier891Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.989597,exponentBits,mantissaBits-1));
        SIGNAL Multiplier892Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.577708,exponentBits,mantissaBits-1));
        SIGNAL Multiplier893Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.618274,exponentBits,mantissaBits-1));
        SIGNAL Multiplier895Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.735141,exponentBits,mantissaBits-1));
        SIGNAL Multiplier896Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.495915,exponentBits,mantissaBits-1));
        SIGNAL Multiplier897Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.993928,exponentBits,mantissaBits-1));
        SIGNAL Multiplier899Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.551341,exponentBits,mantissaBits-1));
        SIGNAL Multiplier900Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.926235,exponentBits,mantissaBits-1));
        SIGNAL Multiplier901Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.616494,exponentBits,mantissaBits-1));
        SIGNAL Multiplier902Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.989597,exponentBits,mantissaBits-1));
        SIGNAL Multiplier903Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.986786,exponentBits,mantissaBits-1));
        SIGNAL Multiplier904Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.464416,exponentBits,mantissaBits-1));
        SIGNAL Multiplier906Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.938375,exponentBits,mantissaBits-1));
        SIGNAL Multiplier908Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.978422,exponentBits,mantissaBits-1));
        SIGNAL Multiplier910Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.773183,exponentBits,mantissaBits-1));
        SIGNAL Multiplier911Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.848299,exponentBits,mantissaBits-1));
        SIGNAL Multiplier912Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.562709,exponentBits,mantissaBits-1));
        SIGNAL Multiplier913Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.988453,exponentBits,mantissaBits-1));
        SIGNAL Multiplier915Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870697,exponentBits,mantissaBits-1));
        SIGNAL Multiplier916Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.945793,exponentBits,mantissaBits-1));
        SIGNAL Multiplier917Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.729204,exponentBits,mantissaBits-1));
        SIGNAL Multiplier918Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870404,exponentBits,mantissaBits-1));
        SIGNAL Multiplier919Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.780732,exponentBits,mantissaBits-1));
        SIGNAL Multiplier920Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.917308,exponentBits,mantissaBits-1));
        SIGNAL Multiplier922Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.631626,exponentBits,mantissaBits-1));
        SIGNAL Multiplier923Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.453222,exponentBits,mantissaBits-1));
        SIGNAL Multiplier924Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.996146,exponentBits,mantissaBits-1));
        SIGNAL Multiplier926Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870697,exponentBits,mantissaBits-1));
        SIGNAL Multiplier927Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.75369,exponentBits,mantissaBits-1));
        SIGNAL Multiplier928Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.936763,exponentBits,mantissaBits-1));
        SIGNAL Multiplier929Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870404,exponentBits,mantissaBits-1));
        SIGNAL Multiplier930Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.933776,exponentBits,mantissaBits-1));
        SIGNAL Multiplier931Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.973389,exponentBits,mantissaBits-1));
        SIGNAL Multiplier933Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.912549,exponentBits,mantissaBits-1));
        SIGNAL Multiplier935Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.973991,exponentBits,mantissaBits-1));
        SIGNAL Multiplier936Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.890735,exponentBits,mantissaBits-1));
        SIGNAL Multiplier937Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.382644,exponentBits,mantissaBits-1));
        SIGNAL Multiplier938Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.998354,exponentBits,mantissaBits-1));
        SIGNAL Multiplier940Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.551341,exponentBits,mantissaBits-1));
        SIGNAL Multiplier941Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.795357,exponentBits,mantissaBits-1));
        SIGNAL Multiplier942Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.948695,exponentBits,mantissaBits-1));
        SIGNAL Multiplier943Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.989597,exponentBits,mantissaBits-1));
        SIGNAL Multiplier944Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.577708,exponentBits,mantissaBits-1));
        SIGNAL Multiplier945Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.98124,exponentBits,mantissaBits-1));
        SIGNAL Multiplier947Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.712179,exponentBits,mantissaBits-1));
        SIGNAL Multiplier948Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.336149,exponentBits,mantissaBits-1));
        SIGNAL Multiplier949Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.99914,exponentBits,mantissaBits-1));
        SIGNAL Multiplier951Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.551341,exponentBits,mantissaBits-1));
        SIGNAL Multiplier952Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.926235,exponentBits,mantissaBits-1));
        SIGNAL Multiplier953Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.981519,exponentBits,mantissaBits-1));
        SIGNAL Multiplier954Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.989597,exponentBits,mantissaBits-1));
        SIGNAL Multiplier955Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.986786,exponentBits,mantissaBits-1));
        SIGNAL Multiplier956Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.995641,exponentBits,mantissaBits-1));
        SIGNAL Multiplier958Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.97267,exponentBits,mantissaBits-1));
        SIGNAL Multiplier960Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.991382,exponentBits,mantissaBits-1));
        SIGNAL Multiplier962Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.56908,exponentBits,mantissaBits-1));
        SIGNAL Multiplier964Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.965849,exponentBits,mantissaBits-1));
        SIGNAL Multiplier965Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.692695,exponentBits,mantissaBits-1));
        SIGNAL Multiplier967Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.880399,exponentBits,mantissaBits-1));
        SIGNAL Multiplier968Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.997554,exponentBits,mantissaBits-1));
        SIGNAL Multiplier969Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.414069,exponentBits,mantissaBits-1));
        SIGNAL Multiplier971Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.91966,exponentBits,mantissaBits-1));
        SIGNAL Multiplier972Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.806938,exponentBits,mantissaBits-1));
        SIGNAL Multiplier974Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.860235,exponentBits,mantissaBits-1));
        SIGNAL Multiplier975Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.989739,exponentBits,mantissaBits-1));
        SIGNAL Multiplier976Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.549861,exponentBits,mantissaBits-1));
        SIGNAL Multiplier979Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.984104,exponentBits,mantissaBits-1));
        SIGNAL Multiplier980Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.793165,exponentBits,mantissaBits-1));
        SIGNAL Multiplier981Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.927417,exponentBits,mantissaBits-1));
        SIGNAL Multiplier983Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.726095,exponentBits,mantissaBits-1));
        SIGNAL Multiplier984Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.98888,exponentBits,mantissaBits-1));
        SIGNAL Multiplier985Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.558577,exponentBits,mantissaBits-1));
        SIGNAL Multiplier987Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.649155,exponentBits,mantissaBits-1));
        SIGNAL Multiplier988Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.975801,exponentBits,mantissaBits-1));
        SIGNAL Multiplier990Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.955917,exponentBits,mantissaBits-1));
        SIGNAL Multiplier991Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.985013,exponentBits,mantissaBits-1));
        SIGNAL Multiplier992Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.592017,exponentBits,mantissaBits-1));
        SIGNAL Multiplier995Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.598812,exponentBits,mantissaBits-1));
        SIGNAL Multiplier997Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.927615,exponentBits,mantissaBits-1));
        SIGNAL Multiplier998Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.792795,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1000Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.907425,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1001Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.948402,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1002Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.83894,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1003Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.898142,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1005Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.826105,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1006Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.838083,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1008Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.965849,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1009Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.692695,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1011Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.880399,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1012Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.997554,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1013Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.414069,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1015Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.91966,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1016Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.806938,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1018Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.860235,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1019Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.989739,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1020Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.549861,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1023Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.932937,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1024Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.793165,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1025Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.927417,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1027Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.726095,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1028Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.98888,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1029Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.558577,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1031Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.649155,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1032Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.975801,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1034Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.955917,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1035Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.985013,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1036Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.592017,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1039Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.782438,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1041Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.750079,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1042Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.947231,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1044Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.907425,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1045Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.74707,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1046Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.617466,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1047Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.981367,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1049Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.826105,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1050Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.898792,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1053Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.914453,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1054Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.965849,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1055Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.692695,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1057Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.880399,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1058Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.966381,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1059Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.690672,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1061Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.91966,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1062Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.806938,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1064Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.860235,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1065Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.94187,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1066Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.763101,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1069Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.924413,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1070Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.793165,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1071Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.927417,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1073Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.726095,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1074Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.909585,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1075Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.82292,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1077Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.649155,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1078Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.975801,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1080Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.955917,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1081Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.790147,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1082Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.929014,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1085Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.798666,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1087Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.927615,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1088Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.792795,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1090Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.807766,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1091Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.907576,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1092Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.83894,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1093Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.898142,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1095Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.919167,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1096Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.781132,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1098Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.965849,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1099Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.692695,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1101Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.880399,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1102Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.966381,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1103Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.690672,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1105Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.91966,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1106Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.806938,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1108Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.860235,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1109Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.94187,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1110Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.763101,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1113Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.693688,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1114Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.793165,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1115Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.927417,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1117Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.726095,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1118Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.909585,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1119Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.82292,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1121Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.649155,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1122Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.975801,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1124Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.955917,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1125Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.790147,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1126Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.929014,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1129Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.965586,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1131Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.750079,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1132Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.947231,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1134Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.807766,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1135Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.825885,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1136Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.617466,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1137Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.981367,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1139Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.919167,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1140Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.93358,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1143Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.815442,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1147Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.848299,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1148Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.895308,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1149Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.842608,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1151Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870697,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1152Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.945793,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1153Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.95487,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1154Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870404,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1155Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.780732,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1156Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.810846,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1158Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.991361,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1159Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.669241,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1160Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.97158,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1162Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870697,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1163Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.75369,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1164Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.77448,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1165Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870404,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1166Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.933776,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1167Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.660973,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1169Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870239,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1171Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.94472,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1172Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.890735,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1173Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.689002,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1174Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.966814,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1176Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.551341,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1177Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.795357,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1178Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.746308,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1179Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.989597,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1180Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.577708,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1181Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.618274,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1183Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.952809,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1184Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.495915,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1185Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.993928,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1187Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.551341,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1188Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.926235,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1189Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.616494,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1190Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.989597,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1191Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.986786,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1192Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.464416,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1194Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.770987,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1196Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.827729,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1198Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.579175,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1199Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.848299,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1200Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.562709,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1201Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.988453,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1203Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870697,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1204Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.945793,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1205Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.729204,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1206Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870404,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1207Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.780732,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1208Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.917308,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1210Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.979033,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1211Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.453222,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1212Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.996146,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1214Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870697,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1215Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.75369,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1216Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.936763,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1217Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870404,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1218Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.933776,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1219Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.973389,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1221Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.818419,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1223Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.766253,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1224Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.890735,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1225Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.382644,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1226Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.998354,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1228Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.551341,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1229Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.795357,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1230Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.948695,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1231Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.989597,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1232Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.577708,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1233Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.98124,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1235Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.960334,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1236Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.336149,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1237Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.99914,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1239Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.551341,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1240Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.926235,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1241Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.981519,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1242Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.989597,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1243Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.986786,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1244Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.995641,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1246Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.664315,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1248Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.634118,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1250Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.760169,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1252Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.970921,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1253Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.67214,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1255Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.98927,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1256Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.997554,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1257Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.414069,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1259Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.853307,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1260Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.886527,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1262Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.554692,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1263Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.989739,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1264Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.549861,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1267Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.994862,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1268Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.817897,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1269Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.912886,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1271Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.976301,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1272Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.98888,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1273Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.558577,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1275Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.731617,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1276Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.954043,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1278Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.646579,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1279Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.985013,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1280Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.592017,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1283Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.479802,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1285Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.807423,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1286Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.919372,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1288Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.694473,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1289Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.843444,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1290Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.682797,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1291Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.968381,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1293Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.965376,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1294Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.697447,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1296Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.970921,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1297Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.67214,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1299Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.98927,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1300Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.997554,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1301Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.414069,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1303Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.853307,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1304Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.886527,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1306Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.554692,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1307Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.989739,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1308Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.549861,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1311Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.970629,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1312Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.817897,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1313Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.912886,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1315Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.976301,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1316Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.98888,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1317Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.558577,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1319Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.731617,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1320Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.954043,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1322Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.646579,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1323Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.985013,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1324Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.592017,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1327Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.673404,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1329Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.62336,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1330Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.980424,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1332Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.694473,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1333Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.894649,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1334Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.482891,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1335Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.994693,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1337Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.965376,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1338Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.964572,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1341Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.952231,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1342Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.970921,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1343Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.67214,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1345Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.98927,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1346Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.966381,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1347Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.690672,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1349Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.853307,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1350Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.886527,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1352Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.554692,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1353Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.94187,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1354Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.763101,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1357Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.951966,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1358Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.817897,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1359Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.912886,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1361Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.976301,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1362Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.909585,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1363Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.82292,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1365Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.731617,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1366Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.954043,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1368Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.646579,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1369Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.790147,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1370Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.929014,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1373Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.7375,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1375Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.807423,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1376Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.919372,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1378Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.579487,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1379Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.790558,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1380Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.682797,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1381Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.968381,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1383Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.986575,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1384Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.578242,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1386Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.970921,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1387Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.67214,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1389Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.98927,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1390Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.966381,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1391Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.690672,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1393Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.853307,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1394Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.886527,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1396Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.554692,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1397Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.94187,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1398Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.763101,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1401Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.840616,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1402Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.817897,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1403Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.912886,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1405Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.976301,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1406Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.909585,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1407Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.82292,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1409Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.731617,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1410Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.954043,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1412Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.646579,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1413Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.790147,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1414Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.929014,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1417Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.896858,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1419Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.62336,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1420Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.980424,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1422Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.579487,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1423Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.928799,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1424Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.482891,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1425Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.994693,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1427Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.986575,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1428Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.986723,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1431Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.736765,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1433Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.848299,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1434Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.895308,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1435Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.842608,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1437Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870697,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1438Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.945793,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1439Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.95487,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1440Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870404,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1441Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.780732,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1442Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.810846,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1444Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.991361,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1445Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.669241,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1446Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.97158,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1448Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870697,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1449Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.75369,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1450Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.77448,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1451Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870404,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1452Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.933776,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1453Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.660973,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1455Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870239,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1457Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.756327,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1458Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.890735,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1459Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.689002,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1460Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.966814,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1462Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.551341,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1463Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.795357,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1464Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.746308,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1465Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.989597,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1466Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.577708,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1467Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.618274,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1469Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.952809,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1470Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.495915,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1471Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.993928,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1473Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.551341,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1474Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.926235,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1475Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.616494,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1476Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.989597,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1477Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.986786,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1478Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.464416,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1480Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.770987,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1482Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.906302,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1484Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.923601,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1485Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.848299,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1486Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.562709,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1487Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.988453,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1489Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870697,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1490Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.945793,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1491Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.729204,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1492Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870404,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1493Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.780732,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1494Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.917308,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1496Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.979033,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1497Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.453222,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1498Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.996146,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1500Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870697,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1501Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.75369,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1502Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.936763,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1503Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870404,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1504Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.933776,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1505Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.973389,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1507Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.818419,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1509Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.940496,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1510Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.890735,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1511Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.382644,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1512Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.998354,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1514Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.551341,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1515Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.795357,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1516Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.948695,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1517Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.989597,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1518Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.577708,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1519Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.98124,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1521Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.960334,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1522Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.336149,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1523Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.99914,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1525Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.551341,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1526Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.926235,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1527Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.981519,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1528Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.989597,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1529Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.986786,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1530Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.995641,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1532Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.664315,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1534Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.978597,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1536Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.974456,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1538Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.970921,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1539Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.67214,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1541Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.98927,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1542Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.997554,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1543Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.414069,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1545Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.853307,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1546Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.886527,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1548Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.554692,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1549Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.989739,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1550Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.549861,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1553Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.994862,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1554Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.817897,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1555Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.912886,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1557Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.976301,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1558Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.98888,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1559Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.558577,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1561Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.731617,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1562Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.954043,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1564Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.646579,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1565Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.985013,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1566Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.592017,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1569Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.479802,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1571Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.807423,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1572Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.919372,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1574Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.694473,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1575Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.843444,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1576Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.682797,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1577Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.968381,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1579Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.965376,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1580Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.697447,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1582Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.970921,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1583Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.67214,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1585Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.98927,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1586Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.997554,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1587Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.414069,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1589Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.853307,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1590Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.886527,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1592Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.554692,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1593Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.989739,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1594Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.549861,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1597Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.970629,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1598Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.817897,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1599Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.912886,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1601Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.976301,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1602Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.98888,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1603Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.558577,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1605Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.731617,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1606Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.954043,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1608Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.646579,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1609Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.985013,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1610Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.592017,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1613Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.673404,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1615Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.62336,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1616Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.980424,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1618Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.694473,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1619Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.894649,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1620Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.482891,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1621Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.994693,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1623Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.965376,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1624Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.964572,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1627Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.768486,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1628Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.970921,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1629Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.67214,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1631Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.98927,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1632Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.966381,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1633Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.690672,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1635Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.853307,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1636Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.886527,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1638Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.554692,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1639Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.94187,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1640Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.763101,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1643Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.951966,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1644Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.817897,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1645Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.912886,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1647Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.976301,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1648Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.909585,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1649Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.82292,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1651Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.731617,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1652Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.954043,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1654Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.646579,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1655Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.790147,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1656Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.929014,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1659Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.7375,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1661Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.807423,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1662Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.919372,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1664Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.579487,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1665Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.790558,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1666Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.682797,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1667Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.968381,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1669Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.986575,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1670Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.578242,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1672Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.970921,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1673Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.67214,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1675Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.98927,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1676Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.966381,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1677Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.690672,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1679Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.853307,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1680Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.886527,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1682Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.554692,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1683Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.94187,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1684Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.763101,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1687Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.840616,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1688Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.817897,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1689Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.912886,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1691Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.976301,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1692Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.909585,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1693Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.82292,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1695Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.731617,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1696Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.954043,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1698Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.646579,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1699Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.790147,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1700Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.929014,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1703Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.896858,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1705Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.62336,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1706Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.980424,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1708Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.579487,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1709Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.928799,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1710Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.482891,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1711Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.994693,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1713Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.986575,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1714Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.986723,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1717Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.939505,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1720Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.848299,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1721Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.895308,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1722Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.842608,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1724Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870697,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1725Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.945793,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1726Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.95487,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1727Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870404,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1728Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.780732,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1729Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.810846,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1731Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.531606,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1732Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.669241,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1733Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.97158,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1735Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870697,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1736Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.75369,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1737Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.77448,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1738Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870404,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1739Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.933776,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1740Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.660973,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1742Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870862,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1744Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.85073,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1745Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.890735,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1746Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.689002,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1747Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.966814,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1749Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.551341,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1750Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.795357,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1751Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.746308,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1752Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.989597,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1753Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.577708,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1754Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.618274,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1756Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.735141,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1757Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.495915,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1758Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.993928,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1760Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.551341,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1761Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.926235,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1762Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.616494,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1763Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.989597,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1764Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.986786,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1765Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.464416,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1767Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.938375,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1769Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.635106,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1771Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.677835,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1772Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.848299,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1773Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.562709,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1774Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.988453,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1776Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870697,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1777Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.945793,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1778Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.729204,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1779Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870404,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1780Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.780732,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1781Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.917308,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1783Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.631626,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1784Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.453222,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1785Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.996146,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1787Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870697,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1788Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.75369,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1789Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.936763,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1790Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870404,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1791Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.933776,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1792Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.973389,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1794Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.912549,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1796Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.658116,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1797Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.890735,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1798Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.382644,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1799Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.998354,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1801Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.551341,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1802Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.795357,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1803Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.948695,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1804Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.989597,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1805Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.577708,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1806Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.98124,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1808Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.712179,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1809Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.336149,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1810Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.99914,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1812Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.551341,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1813Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.926235,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1814Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.981519,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1815Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.989597,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1816Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.986786,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1817Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.995641,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1819Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.97267,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1821Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.53135,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1823Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.816772,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1825Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.965849,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1826Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.692695,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1828Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.880399,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1829Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.997554,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1830Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.414069,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1832Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.91966,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1833Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.806938,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1835Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.860235,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1836Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.989739,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1837Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.549861,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1840Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.984104,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1841Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.793165,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1842Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.927417,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1844Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.726095,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1845Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.98888,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1846Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.558577,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1848Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.649155,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1849Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.975801,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1851Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.955917,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1852Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.985013,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1853Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.592017,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1856Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.598812,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1858Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.807423,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1859Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.919372,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1861Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.694473,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1862Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.843444,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1863Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.682797,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1864Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.968381,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1866Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.965376,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1867Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.697447,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1869Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.965849,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1870Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.692695,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1872Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.880399,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1873Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.997554,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1874Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.414069,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1876Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.91966,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1877Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.806938,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1879Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.860235,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1880Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.989739,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1881Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.549861,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1884Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.932937,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1885Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.793165,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1886Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.927417,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1888Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.726095,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1889Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.98888,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1890Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.558577,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1892Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.649155,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1893Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.975801,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1895Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.955917,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1896Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.985013,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1897Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.592017,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1900Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.782438,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1902Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.62336,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1903Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.980424,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1905Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.694473,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1906Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.894649,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1907Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.482891,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1908Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.994693,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1910Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.965376,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1911Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.964572,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1914Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.926565,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1915Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.965849,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1916Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.692695,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1918Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.880399,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1919Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.966381,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1920Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.690672,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1922Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.91966,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1923Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.806938,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1925Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.860235,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1926Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.94187,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1927Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.763101,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1930Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.924413,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1931Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.793165,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1932Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.927417,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1934Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.726095,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1935Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.909585,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1936Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.82292,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1938Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.649155,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1939Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.975801,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1941Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.955917,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1942Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.790147,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1943Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.929014,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1946Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.798666,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1948Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.807423,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1949Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.919372,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1951Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.579487,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1952Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.790558,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1953Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.682797,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1954Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.968381,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1956Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.986575,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1957Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.578242,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1959Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.965849,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1960Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.692695,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1962Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.880399,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1963Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.966381,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1964Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.690672,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1966Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.91966,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1967Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.806938,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1969Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.860235,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1970Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.94187,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1971Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.763101,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1974Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.693688,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1975Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.793165,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1976Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.927417,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1978Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.726095,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1979Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.909585,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1980Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.82292,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1982Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.649155,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1983Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.975801,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1985Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.955917,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1986Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.790147,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1987Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.929014,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1990Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.965586,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1992Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.62336,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1993Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.980424,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1995Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.579487,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1996Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.928799,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1997Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.482891,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1998Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.994693,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2000Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.986575,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2001Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.986723,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2004Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.794749,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2006Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.848299,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2007Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.895308,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2008Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.842608,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2010Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870697,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2011Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.945793,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2012Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.95487,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2013Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870404,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2014Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.780732,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2015Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.810846,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2017Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.531606,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2018Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.669241,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2019Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.97158,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2021Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870697,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2022Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.75369,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2023Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.77448,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2024Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870404,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2025Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.933776,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2026Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.660973,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2028Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870862,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2030Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.888715,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2031Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.890735,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2032Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.689002,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2033Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.966814,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2035Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.551341,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2036Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.795357,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2037Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.746308,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2038Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.989597,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2039Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.577708,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2040Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.618274,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2042Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.735141,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2043Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.495915,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2044Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.993928,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2046Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.551341,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2047Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.926235,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2048Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.616494,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2049Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.989597,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2050Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.986786,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2051Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.464416,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2053Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.938375,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2055Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.978422,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2057Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.937366,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2058Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.848299,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2059Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.562709,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2060Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.988453,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2062Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870697,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2063Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.945793,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2064Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.729204,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2065Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870404,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2066Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.780732,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2067Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.917308,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2069Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.631626,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2070Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.453222,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2071Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.996146,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2073Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870697,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2074Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.75369,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2075Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.936763,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2076Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.870404,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2077Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.933776,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2078Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.973389,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2080Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.912549,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2082Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.973991,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2083Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.890735,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2084Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.382644,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2085Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.998354,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2087Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.551341,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2088Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.795357,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2089Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.948695,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2090Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.989597,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2091Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.577708,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2092Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.98124,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2094Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.712179,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2095Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.336149,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2096Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.99914,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2098Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.551341,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2099Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.926235,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2100Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.981519,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2101Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.989597,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2102Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.986786,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2103Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.995641,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2105Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.97267,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2107Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.991382,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2109Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.987767,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2111Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.965849,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2112Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.692695,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2114Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.880399,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2115Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.997554,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2116Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.414069,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2118Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.91966,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2119Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.806938,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2121Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.860235,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2122Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.989739,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2123Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.549861,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2126Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.984104,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2127Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.793165,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2128Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.927417,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2130Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.726095,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2131Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.98888,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2132Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.558577,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2134Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.649155,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2135Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.975801,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2137Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.955917,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2138Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.985013,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2139Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.592017,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2142Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.598812,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2144Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.807423,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2145Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.919372,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2147Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.694473,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2148Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.843444,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2149Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.682797,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2150Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.968381,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2152Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.965376,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2153Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.697447,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2155Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.965849,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2156Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.692695,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2158Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.880399,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2159Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.997554,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2160Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.414069,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2162Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.91966,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2163Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.806938,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2165Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.860235,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2166Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.989739,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2167Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.549861,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2170Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.932937,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2171Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.793165,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2172Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.927417,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2174Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.726095,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2175Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.98888,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2176Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.558577,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2178Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.649155,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2179Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.975801,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2181Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.955917,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2182Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.985013,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2183Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.592017,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2186Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.782438,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2188Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.62336,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2189Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.980424,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2191Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.694473,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2192Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.894649,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2193Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.482891,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2194Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.994693,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2196Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.965376,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2197Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.964572,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2200Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.625034,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2201Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.965849,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2202Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.692695,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2204Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.880399,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2205Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.966381,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2206Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.690672,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2208Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.91966,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2209Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.806938,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2211Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.860235,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2212Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.94187,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2213Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.763101,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2216Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.924413,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2217Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.793165,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2218Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.927417,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2220Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.726095,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2221Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.909585,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2222Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.82292,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2224Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.649155,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2225Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.975801,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2227Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.955917,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2228Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.790147,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2229Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.929014,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2232Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.798666,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2234Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.807423,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2235Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.919372,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2237Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.579487,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2238Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.790558,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2239Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.682797,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2240Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.968381,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2242Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.986575,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2243Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.578242,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2245Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.965849,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2246Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.692695,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2248Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.880399,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2249Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.966381,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2250Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.690672,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2252Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.91966,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2253Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.806938,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2255Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.860235,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2256Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.94187,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2257Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.763101,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2260Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.693688,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2261Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.793165,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2262Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.927417,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2264Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.726095,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2265Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.909585,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2266Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.82292,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2268Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.649155,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2269Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.975801,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2271Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.955917,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2272Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.790147,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2273Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.929014,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2276Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.965586,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2278Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.62336,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2279Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.980424,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2281Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.579487,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2282Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.928799,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2283Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.482891,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2284Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.994693,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2286Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.986575,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2287Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.986723,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2290Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.980149,exponentBits,mantissaBits-1));
        
BEGIN
    PROCESS (clk,rst) IS
    BEGIN 
        IF rst = '1' THEN
    mbRightSHR2293_2955Input <= (others=>'0');
            mbRightSHR1146_1477Input <= (others=>'0');
mbRightSHR2292_2953Input <= (others=>'0');
            mbRightSHR1719_2215Input <= (others=>'0');
            mbRightSHR1145_1475Input <= (others=>'0');
            mbRightSHR572_737Input <= (others=>'0');
mbRightSHR2110_2711Input <= (others=>'0');
            mbRightSHR1824_2343Input <= (others=>'0');
            mbRightSHR1537_1973Input <= (others=>'0');
            mbRightSHR1251_1605Input <= (others=>'0');
            mbRightSHR963_1233Input <= (others=>'0');
            mbRightSHR677_865Input <= (others=>'0');
            mbRightSHR390_495Input <= (others=>'0');
            mbRightSHR104_127Input <= (others=>'0');
mbRightSHR2003_2580Input <= (others=>'0');
            mbRightSHR1913_2461Input <= (others=>'0');
            mbRightSHR1430_1842Input <= (others=>'0');
            mbRightSHR1340_1723Input <= (others=>'0');
            mbRightSHR856_1102Input <= (others=>'0');
            mbRightSHR766_983Input <= (others=>'0');
            mbRightSHR283_364Input <= (others=>'0');
            mbRightSHR193_245Input <= (others=>'0');
mbRightSHR961_1230Input <= (others=>'0');
            mbRightSHR909_1167Input <= (others=>'0');
            mbRightSHR675_862Input <= (others=>'0');
            mbRightSHR623_799Input <= (others=>'0');
            mbRightSHR388_492Input <= (others=>'0');
            mbRightSHR336_429Input <= (others=>'0');
            mbRightSHR102_124Input <= (others=>'0');
            mbRightSHR50_61Input <= (others=>'0');
mbRightSHR844_1086Input <= (others=>'0');
            mbRightSHR800_1028Input <= (others=>'0');
            mbRightSHR754_967Input <= (others=>'0');
            mbRightSHR710_909Input <= (others=>'0');
            mbRightSHR271_348Input <= (others=>'0');
            mbRightSHR227_290Input <= (others=>'0');
            mbRightSHR181_229Input <= (others=>'0');
            mbRightSHR137_171Input <= (others=>'0');
mbRightSHR25_Input2_30Input <= (others=>'0');
            mbRightSHR0_Input2_0Input <= (others=>'0');
mbRightSHR1336_1717Input <= (others=>'0');
            mbRightSHR1331_1711Input <= (others=>'0');
            mbRightSHR798_1025Input <= (others=>'0');
            mbRightSHR782_1004Input <= (others=>'0');
            mbRightSHR1292_1659Input <= (others=>'0');
            mbRightSHR1287_1653Input <= (others=>'0');
            mbRightSHR708_906Input <= (others=>'0');
            mbRightSHR692_885Input <= (others=>'0');
            mbRightSHR225_287Input <= (others=>'0');
            mbRightSHR209_266Input <= (others=>'0');
            mbRightSHR135_168Input <= (others=>'0');
            mbRightSHR119_147Input <= (others=>'0');
            mbRightSHR189_239Input <= (others=>'0');
            mbRightSHR184_233Input <= (others=>'0');
            mbRightSHR145_181Input <= (others=>'0');
            mbRightSHR140_175Input <= (others=>'0');
mbRightSHR1335_Input2_1715Input <= (others=>'0');
            mbRightSHR1334_Input2_1714Input <= (others=>'0');
            mbRightSHR1330_Input2_1709Input <= (others=>'0');
            mbRightSHR1329_Input2_1708Input <= (others=>'0');
            mbRightSHR1291_Input2_1657Input <= (others=>'0');
            mbRightSHR1290_Input2_1656Input <= (others=>'0');
            mbRightSHR1286_Input2_1651Input <= (others=>'0');
            mbRightSHR1285_Input2_1650Input <= (others=>'0');
            mbRightSHR91_110Input <= (others=>'0');
            mbRightSHR80_97Input <= (others=>'0');
            mbRightSHR66_80Input <= (others=>'0');
            mbRightSHR55_67Input <= (others=>'0');
            mbRightSHR39_47Input <= (others=>'0');
            mbRightSHR28_34Input <= (others=>'0');
            mbRightSHR14_17Input <= (others=>'0');
            mbRightSHR3_4Input <= (others=>'0');
            mbRightSHR188_Input2_237Input <= (others=>'0');
            mbRightSHR187_Input2_236Input <= (others=>'0');
            mbRightSHR183_Input2_231Input <= (others=>'0');
            mbRightSHR182_Input2_230Input <= (others=>'0');
            mbRightSHR144_Input2_179Input <= (others=>'0');
            mbRightSHR143_Input2_178Input <= (others=>'0');
            mbRightSHR139_Input2_173Input <= (others=>'0');
            mbRightSHR138_Input2_172Input <= (others=>'0');
mbRightSHR223_Input2_283Input <= (others=>'0');
            mbRightSHR222_Input2_282Input <= (others=>'0');
            mbRightSHR703_899Input <= (others=>'0');
            mbRightSHR216_Input2_274Input <= (others=>'0');
            mbRightSHR215_Input2_273Input <= (others=>'0');
            mbRightSHR696_890Input <= (others=>'0');
            mbRightSHR207_Input2_262Input <= (others=>'0');
            mbRightSHR206_Input2_261Input <= (others=>'0');
            mbRightSHR687_878Input <= (others=>'0');
            mbRightSHR200_Input2_253Input <= (others=>'0');
            mbRightSHR199_Input2_252Input <= (others=>'0');
            mbRightSHR680_869Input <= (others=>'0');
            mbRightSHR133_Input2_164Input <= (others=>'0');
            mbRightSHR132_Input2_163Input <= (others=>'0');
            mbRightSHR126_Input2_155Input <= (others=>'0');
            mbRightSHR125_Input2_154Input <= (others=>'0');
            mbRightSHR117_Input2_143Input <= (others=>'0');
            mbRightSHR116_Input2_142Input <= (others=>'0');
            mbRightSHR110_Input2_134Input <= (others=>'0');
            mbRightSHR109_Input2_133Input <= (others=>'0');
            mbRightSHR90_Input2_108Input <= (others=>'0');
            mbRightSHR89_Input2_107Input <= (others=>'0');
            mbRightSHR79_Input2_95Input <= (others=>'0');
            mbRightSHR78_Input2_94Input <= (others=>'0');
            mbRightSHR65_Input2_78Input <= (others=>'0');
            mbRightSHR64_Input2_77Input <= (others=>'0');
            mbRightSHR54_Input2_65Input <= (others=>'0');
            mbRightSHR53_Input2_64Input <= (others=>'0');
            mbRightSHR38_Input2_45Input <= (others=>'0');
            mbRightSHR37_Input2_44Input <= (others=>'0');
            mbRightSHR27_Input2_32Input <= (others=>'0');
            mbRightSHR26_Input2_31Input <= (others=>'0');
            mbRightSHR13_Input2_15Input <= (others=>'0');
            mbRightSHR12_Input2_14Input <= (others=>'0');
            mbRightSHR2_Input2_2Input <= (others=>'0');
            mbRightSHR1_Input2_1Input <= (others=>'0');
            mbRightSHR130_161Input <= (others=>'0');
            mbRightSHR123_152Input <= (others=>'0');
            mbRightSHR114_140Input <= (others=>'0');
            mbRightSHR107_131Input <= (others=>'0');
mbRightSHR32_Input2_38Input <= (others=>'0');
            mbRightSHR29_Input2_35Input <= (others=>'0');
            mbRightSHR7_Input2_8Input <= (others=>'0');
            mbRightSHR4_Input2_5Input <= (others=>'0');
mb_D_FFMultiplier21_702_0Input <= (others=>'0');
            mb_D_FFMultiplier21_701_0Input <= (others=>'0');
            mb_D_FFMultiplier21_695_0Input <= (others=>'0');
            mb_D_FFMultiplier21_694_0Input <= (others=>'0');
            mb_D_FFMultiplier21_686_0Input <= (others=>'0');
            mb_D_FFMultiplier21_685_0Input <= (others=>'0');
            mb_D_FFMultiplier21_679_0Input <= (others=>'0');
            mb_D_FFMultiplier21_678_0Input <= (others=>'0');
            mb_D_FFMultiplier21_129_0Input <= (others=>'0');
            mb_D_FFMultiplier21_128_0Input <= (others=>'0');
            mb_D_FFMultiplier21_122_0Input <= (others=>'0');
            mb_D_FFMultiplier21_121_0Input <= (others=>'0');
            mb_D_FFMultiplier21_113_0Input <= (others=>'0');
            mb_D_FFMultiplier21_112_0Input <= (others=>'0');
            mb_D_FFMultiplier21_106_0Input <= (others=>'0');
            mb_D_FFMultiplier21_105_0Input <= (others=>'0');
        ELSIF rising_edge(clk) and rst = '0' and enable = '1' THEN
            mbRightSHR2293_2955Input <= vb14;
            mbRightSHR1146_1477Input <= v14;
mbRightSHR2292_2953Input <= vb6;
            mbRightSHR1719_2215Input <= v6;
            mbRightSHR1145_1475Input <= vb6;
            mbRightSHR572_737Input <= v6;
mbRightSHR2110_2711Input <= vb16;
            mbRightSHR1824_2343Input <= v16;
            mbRightSHR1537_1973Input <= vb16;
            mbRightSHR1251_1605Input <= v16;
            mbRightSHR963_1233Input <= vb16;
            mbRightSHR677_865Input <= v16;
            mbRightSHR390_495Input <= vb16;
            mbRightSHR104_127Input <= v16;
mbRightSHR2003_2580Input <= vb15;
            mbRightSHR1913_2461Input <= v15;
            mbRightSHR1430_1842Input <= vb15;
            mbRightSHR1340_1723Input <= v15;
            mbRightSHR856_1102Input <= vb15;
            mbRightSHR766_983Input <= v15;
            mbRightSHR283_364Input <= vb15;
            mbRightSHR193_245Input <= v15;
mbRightSHR961_1230Input <= vb5;
            mbRightSHR909_1167Input <= v5;
            mbRightSHR675_862Input <= vb5;
            mbRightSHR623_799Input <= v5;
            mbRightSHR388_492Input <= vb5;
            mbRightSHR336_429Input <= v5;
            mbRightSHR102_124Input <= vb5;
            mbRightSHR50_61Input <= v5;
mbRightSHR844_1086Input <= vb10;
            mbRightSHR800_1028Input <= v10;
            mbRightSHR754_967Input <= vb10;
            mbRightSHR710_909Input <= v10;
            mbRightSHR271_348Input <= vb10;
            mbRightSHR227_290Input <= v10;
            mbRightSHR181_229Input <= vb10;
            mbRightSHR137_171Input <= v10;
mbRightSHR25_Input2_30Input <= vb4;
            mbRightSHR0_Input2_0Input <= v4;
mbRightSHR1336_1717Input <= vb9;
            mbRightSHR1331_1711Input <= v9;
            mbRightSHR798_1025Input <= vb13;
            mbRightSHR782_1004Input <= v13;
            mbRightSHR1292_1659Input <= vb9;
            mbRightSHR1287_1653Input <= v9;
            mbRightSHR708_906Input <= vb13;
            mbRightSHR692_885Input <= v13;
            mbRightSHR225_287Input <= vb13;
            mbRightSHR209_266Input <= v13;
            mbRightSHR135_168Input <= vb13;
            mbRightSHR119_147Input <= v13;
            mbRightSHR189_239Input <= vb9;
            mbRightSHR184_233Input <= v9;
            mbRightSHR145_181Input <= vb9;
            mbRightSHR140_175Input <= v9;
mbRightSHR1335_Input2_1715Input <= vb1;
            mbRightSHR1334_Input2_1714Input <= v1;
            mbRightSHR1330_Input2_1709Input <= vb1;
            mbRightSHR1329_Input2_1708Input <= v1;
            mbRightSHR1291_Input2_1657Input <= vb1;
            mbRightSHR1290_Input2_1656Input <= v1;
            mbRightSHR1286_Input2_1651Input <= vb1;
            mbRightSHR1285_Input2_1650Input <= v1;
            mbRightSHR91_110Input <= vb7;
            mbRightSHR80_97Input <= v7;
            mbRightSHR66_80Input <= vb7;
            mbRightSHR55_67Input <= v7;
            mbRightSHR39_47Input <= vb7;
            mbRightSHR28_34Input <= v7;
            mbRightSHR14_17Input <= vb7;
            mbRightSHR3_4Input <= v7;
            mbRightSHR188_Input2_237Input <= vb1;
            mbRightSHR187_Input2_236Input <= v1;
            mbRightSHR183_Input2_231Input <= vb1;
            mbRightSHR182_Input2_230Input <= v1;
            mbRightSHR144_Input2_179Input <= vb1;
            mbRightSHR143_Input2_178Input <= v1;
            mbRightSHR139_Input2_173Input <= vb1;
            mbRightSHR138_Input2_172Input <= v1;
mbRightSHR223_Input2_283Input <= vb2;
            mbRightSHR222_Input2_282Input <= v2;
            mbRightSHR703_899Input <= vb12;
            mbRightSHR216_Input2_274Input <= vb2;
            mbRightSHR215_Input2_273Input <= v2;
            mbRightSHR696_890Input <= v12;
            mbRightSHR207_Input2_262Input <= vb2;
            mbRightSHR206_Input2_261Input <= v2;
            mbRightSHR687_878Input <= vb12;
            mbRightSHR200_Input2_253Input <= vb2;
            mbRightSHR199_Input2_252Input <= v2;
            mbRightSHR680_869Input <= v12;
            mbRightSHR133_Input2_164Input <= vb2;
            mbRightSHR132_Input2_163Input <= v2;
            mbRightSHR126_Input2_155Input <= vb2;
            mbRightSHR125_Input2_154Input <= v2;
            mbRightSHR117_Input2_143Input <= vb2;
            mbRightSHR116_Input2_142Input <= v2;
            mbRightSHR110_Input2_134Input <= vb2;
            mbRightSHR109_Input2_133Input <= v2;
            mbRightSHR90_Input2_108Input <= vb8;
            mbRightSHR89_Input2_107Input <= v8;
            mbRightSHR79_Input2_95Input <= vb8;
            mbRightSHR78_Input2_94Input <= v8;
            mbRightSHR65_Input2_78Input <= vb8;
            mbRightSHR64_Input2_77Input <= v8;
            mbRightSHR54_Input2_65Input <= vb8;
            mbRightSHR53_Input2_64Input <= v8;
            mbRightSHR38_Input2_45Input <= vb8;
            mbRightSHR37_Input2_44Input <= v8;
            mbRightSHR27_Input2_32Input <= vb8;
            mbRightSHR26_Input2_31Input <= v8;
            mbRightSHR13_Input2_15Input <= vb8;
            mbRightSHR12_Input2_14Input <= v8;
            mbRightSHR2_Input2_2Input <= vb8;
            mbRightSHR1_Input2_1Input <= v8;
            mbRightSHR130_161Input <= vb12;
            mbRightSHR123_152Input <= v12;
            mbRightSHR114_140Input <= vb12;
            mbRightSHR107_131Input <= v12;
mbRightSHR32_Input2_38Input <= vb3;
            mbRightSHR29_Input2_35Input <= v3;
            mbRightSHR7_Input2_8Input <= vb3;
            mbRightSHR4_Input2_5Input <= v3;
mb_D_FFMultiplier21_702_0Input <= vb11;
            mb_D_FFMultiplier21_701_0Input <= v11;
            mb_D_FFMultiplier21_695_0Input <= vb11;
            mb_D_FFMultiplier21_694_0Input <= v11;
            mb_D_FFMultiplier21_686_0Input <= vb11;
            mb_D_FFMultiplier21_685_0Input <= v11;
            mb_D_FFMultiplier21_679_0Input <= vb11;
            mb_D_FFMultiplier21_678_0Input <= v11;
            mb_D_FFMultiplier21_129_0Input <= vb11;
            mb_D_FFMultiplier21_128_0Input <= v11;
            mb_D_FFMultiplier21_122_0Input <= vb11;
            mb_D_FFMultiplier21_121_0Input <= v11;
            mb_D_FFMultiplier21_113_0Input <= vb11;
            mb_D_FFMultiplier21_112_0Input <= v11;
            mb_D_FFMultiplier21_106_0Input <= vb11;
            mb_D_FFMultiplier21_105_0Input <= v11;
        END IF;

    END PROCESS;

    MBRightSHR_Float_0_Input10: entity work.MBRightSHR(rtl)
    GENERIC MAP (89, NumberOfBits)
    PORT MAP (clk, rst, Multiplier0Weight, mbRightSHR0_Input1_0Output);

    MB_D_FF_Float_0_0_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR0_Input1_0Output, Multiplier0WeightOutput);

    InputIEEE_Float_0_0: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier0WeightOutput, flopocoMultiplier0WeightOutput);

    MB_D_FF_Float_0_0_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier0WeightOutput, flopocoMultiplier0WeightInput);

    Multiplier_Float_0: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier0WeightInput, mb_D_FF0_0MultiplierStage2Output, Multiplier0_Output_0);

    MBRightSHR_Float_0_Input2_0: entity work.MBRightSHR(rtl)
    GENERIC MAP (89, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR0_Input2_0Input, mbRightSHR0_Input2_0Output);

    MB_D_FF_Float_0_0_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR0_Input2_0Output, mb_D_FF0_0MultiplierStage1Output);

    MB_D_FF_Float_0_0_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF0_0MultiplierStage1Output, mb_D_FF0_0MultiplierStage2Output);

    MBRightSHR_Float_1_Input11: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits)
    PORT MAP (clk, rst, Multiplier1Weight, mbRightSHR1_Input1_1Output);

    MB_D_FF_Float_1_1_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR1_Input1_1Output, Multiplier1WeightOutput);

    InputIEEE_Float_1_1: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier1WeightOutput, flopocoMultiplier1WeightOutput);

    MB_D_FF_Float_1_1_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier1WeightOutput, flopocoMultiplier1WeightInput);

    Multiplier_Float_1: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier1WeightInput, mb_D_FF1_1MultiplierStage2Output, Multiplier1_Output_1);

    MBRightSHR_Float_1_Input2_1: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR1_Input2_1Input, mbRightSHR1_Input2_1Output);

    MB_D_FF_Float_1_1_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR1_Input2_1Output, mb_D_FF1_1MultiplierStage1Output);

    MB_D_FF_Float_1_1_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1_1MultiplierStage1Output, mb_D_FF1_1MultiplierStage2Output);

    MBRightSHR_Float_2_Input12: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits)
    PORT MAP (clk, rst, Multiplier2Weight, mbRightSHR2_Input1_2Output);

    MB_D_FF_Float_2_2_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR2_Input1_2Output, Multiplier2WeightOutput);

    InputIEEE_Float_2_2: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier2WeightOutput, flopocoMultiplier2WeightOutput);

    MB_D_FF_Float_2_2_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier2WeightOutput, flopocoMultiplier2WeightInput);

    Multiplier_Float_2: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier2WeightInput, mb_D_FF2_2MultiplierStage2Output, Multiplier2_Output_2);

    MBRightSHR_Float_2_Input2_2: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR2_Input2_2Input, mbRightSHR2_Input2_2Output);

    MB_D_FF_Float_2_2_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR2_Input2_2Output, mb_D_FF2_2MultiplierStage1Output);

    MB_D_FF_Float_2_2_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF2_2MultiplierStage1Output, mb_D_FF2_2MultiplierStage2Output);

    MB_D_FF_Float_Adder18_Input1_0_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier2_Output_2, mb_D_FFAdder18_Input1_0_0Output);

    MB_D_FF_Float_0_3_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder18_Input1_0_0Output, mb_D_FF0_3AugendStage1Output);

    MB_D_FF_Float_0_3_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF0_3AugendStage1Output, mb_D_FF0_3AugendStage2Output);

    Adder_Float_0: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF0_3AugendStage2Output, mb_D_FF0_3AddendStage2Output, Adder0_Output_3);

    MB_D_FF_Float_Adder18_Input2_0_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier1_Output_1, mb_D_FFAdder18_Input2_0_0Output);

    MB_D_FF_Float_0_3_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder18_Input2_0_0Output, mb_D_FF0_3AddendStage1Output);

    MB_D_FF_Float_0_3_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF0_3AddendStage1Output, mb_D_FF0_3AddendStage2Output);

    MB_D_FF_Float_Multiplier17_3_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder0_Output_3, mb_D_FFMultiplier17_3_0Output);

    MB_D_FF_Float_3_4_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier17_3_0Output, mb_D_FF3_4MultiplierStage1Output);

    MB_D_FF_Float_3_4_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF3_4MultiplierStage1Output, mb_D_FF3_4MultiplierStage2Output);

    Multiplier_Float_3: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF3_4MultiplierStage2Output, mb_D_FF3_4MultiplicandStage2Output, Multiplier3_Output_4);

    MBRightSHR_Float_3_4: entity work.MBRightSHR(rtl)
    GENERIC MAP (50, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR3_4Input, mbRightSHR3_4Output);

    MB_D_FF_Float_3_4_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR3_4Output, mb_D_FF3_4MultiplicandStage1Output);

    MB_D_FF_Float_3_4_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF3_4MultiplicandStage1Output, mb_D_FF3_4MultiplicandStage2Output);

    MBRightSHR_Float_4_Input15: entity work.MBRightSHR(rtl)
    GENERIC MAP (11, NumberOfBits)
    PORT MAP (clk, rst, Multiplier4Weight, mbRightSHR4_Input1_5Output);

    MB_D_FF_Float_4_5_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR4_Input1_5Output, Multiplier4WeightOutput);

    InputIEEE_Float_4_5: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier4WeightOutput, flopocoMultiplier4WeightOutput);

    MB_D_FF_Float_4_5_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier4WeightOutput, flopocoMultiplier4WeightInput);

    Multiplier_Float_4: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier4WeightInput, mb_D_FF4_5MultiplierStage2Output, Multiplier4_Output_5);

    MBRightSHR_Float_4_Input2_5: entity work.MBRightSHR(rtl)
    GENERIC MAP (11, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR4_Input2_5Input, mbRightSHR4_Input2_5Output);

    MB_D_FF_Float_4_5_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR4_Input2_5Output, mb_D_FF4_5MultiplierStage1Output);

    MB_D_FF_Float_4_5_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF4_5MultiplierStage1Output, mb_D_FF4_5MultiplierStage2Output);

    MB_D_FF_Float_Multiplier19_5_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier4_Output_5, mb_D_FFMultiplier19_5_0Output);

    MB_D_FF_Float_5_6_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier19_5_0Output, mb_D_FF5_6MultiplierStage1Output);

    MB_D_FF_Float_5_6_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF5_6MultiplierStage1Output, mb_D_FF5_6MultiplierStage2Output);

    Multiplier_Float_5: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF5_6MultiplierStage2Output, flopocoMultiplier5WeightInput, Multiplier5_Output_6);

    MBRightSHR_Float_5_6: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits)
    PORT MAP (clk, rst, Multiplier5Weight, mbRightSHR5_6Output);

    MB_D_FF_Float_5_6_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR5_6Output, Multiplier5WeightOutput);

    InputIEEE_Float_5_6: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier5WeightOutput, flopocoMultiplier5WeightOutput);

    MB_D_FF_Float_5_6_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier5WeightOutput, flopocoMultiplier5WeightInput);

    MB_D_FF_Float_Multiplier18_6_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier5_Output_6, mb_D_FFMultiplier18_6_0Output);

    MB_D_FF_Float_6_7_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier18_6_0Output, mb_D_FF6_7MultiplierStage1Output);

    MB_D_FF_Float_6_7_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF6_7MultiplierStage1Output, mb_D_FF6_7MultiplierStage2Output);

    Multiplier_Float_6: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF6_7MultiplierStage2Output, flopocoMultiplier6WeightInput, Multiplier6_Output_7);

    MBRightSHR_Float_6_7: entity work.MBRightSHR(rtl)
    GENERIC MAP (43, NumberOfBits)
    PORT MAP (clk, rst, Multiplier6Weight, mbRightSHR6_7Output);

    MB_D_FF_Float_6_7_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR6_7Output, Multiplier6WeightOutput);

    InputIEEE_Float_6_7: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier6WeightOutput, flopocoMultiplier6WeightOutput);

    MB_D_FF_Float_6_7_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier6WeightOutput, flopocoMultiplier6WeightInput);

    MBRightSHR_Float_7_Input18: entity work.MBRightSHR(rtl)
    GENERIC MAP (11, NumberOfBits)
    PORT MAP (clk, rst, Multiplier7Weight, mbRightSHR7_Input1_8Output);

    MB_D_FF_Float_7_8_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR7_Input1_8Output, Multiplier7WeightOutput);

    InputIEEE_Float_7_8: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier7WeightOutput, flopocoMultiplier7WeightOutput);

    MB_D_FF_Float_7_8_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier7WeightOutput, flopocoMultiplier7WeightInput);

    Multiplier_Float_7: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier7WeightInput, mb_D_FF7_8MultiplierStage2Output, Multiplier7_Output_8);

    MBRightSHR_Float_7_Input2_8: entity work.MBRightSHR(rtl)
    GENERIC MAP (11, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR7_Input2_8Input, mbRightSHR7_Input2_8Output);

    MB_D_FF_Float_7_8_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR7_Input2_8Output, mb_D_FF7_8MultiplierStage1Output);

    MB_D_FF_Float_7_8_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF7_8MultiplierStage1Output, mb_D_FF7_8MultiplierStage2Output);

    MB_D_FF_Float_Multiplier19_8_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier7_Output_8, mb_D_FFMultiplier19_8_0Output);

    MB_D_FF_Float_8_9_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier19_8_0Output, mb_D_FF8_9MultiplierStage1Output);

    MB_D_FF_Float_8_9_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF8_9MultiplierStage1Output, mb_D_FF8_9MultiplierStage2Output);

    Multiplier_Float_8: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF8_9MultiplierStage2Output, flopocoMultiplier8WeightInput, Multiplier8_Output_9);

    MBRightSHR_Float_8_9: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits)
    PORT MAP (clk, rst, Multiplier8Weight, mbRightSHR8_9Output);

    MB_D_FF_Float_8_9_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR8_9Output, Multiplier8WeightOutput);

    InputIEEE_Float_8_9: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier8WeightOutput, flopocoMultiplier8WeightOutput);

    MB_D_FF_Float_8_9_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier8WeightOutput, flopocoMultiplier8WeightInput);

    MB_D_FF_Float_Multiplier18_9_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier8_Output_9, mb_D_FFMultiplier18_9_0Output);

    MB_D_FF_Float_9_10_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier18_9_0Output, mb_D_FF9_10MultiplierStage1Output);

    MB_D_FF_Float_9_10_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF9_10MultiplierStage1Output, mb_D_FF9_10MultiplierStage2Output);

    Multiplier_Float_9: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF9_10MultiplierStage2Output, flopocoMultiplier9WeightInput, Multiplier9_Output_10);

    MBRightSHR_Float_9_10: entity work.MBRightSHR(rtl)
    GENERIC MAP (43, NumberOfBits)
    PORT MAP (clk, rst, Multiplier9Weight, mbRightSHR9_10Output);

    MB_D_FF_Float_9_10_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR9_10Output, Multiplier9WeightOutput);

    InputIEEE_Float_9_10: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier9WeightOutput, flopocoMultiplier9WeightOutput);

    MB_D_FF_Float_9_10_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier9WeightOutput, flopocoMultiplier9WeightInput);

    MB_D_FF_Float_Adder17_Input1_1_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier9_Output_10, mb_D_FFAdder17_Input1_1_0Output);

    MB_D_FF_Float_1_11_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder17_Input1_1_0Output, mb_D_FF1_11AugendStage1Output);

    MB_D_FF_Float_1_11_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1_11AugendStage1Output, mb_D_FF1_11AugendStage2Output);

    Adder_Float_1: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF1_11AugendStage2Output, mb_D_FF1_11AddendStage2Output, Adder1_Output_11);

    MB_D_FF_Float_Adder17_Input2_1_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier6_Output_7, mb_D_FFAdder17_Input2_1_0Output);

    MB_D_FF_Float_1_11_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder17_Input2_1_0Output, mb_D_FF1_11AddendStage1Output);

    MB_D_FF_Float_1_11_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1_11AddendStage1Output, mb_D_FF1_11AddendStage2Output);

    MB_D_FF_Float_Multiplier16_Input1_10_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder1_Output_11, mb_D_FFMultiplier16_Input1_10_0Output);

    MB_D_FF_Float_10_12_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier16_Input1_10_0Output, mb_D_FF10_12MultiplicandStage1Output);

    MB_D_FF_Float_10_12_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF10_12MultiplicandStage1Output, mb_D_FF10_12MultiplicandStage2Output);

    Multiplier_Float_10: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF10_12MultiplicandStage2Output, mb_D_FF10_12MultiplierStage2Output, Multiplier10_Output_12);

    MB_D_FF_Float_Multiplier16_Input2_10_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier3_Output_4, mb_D_FFMultiplier16_Input2_10_0Output);

    MB_D_FF_Float_10_12_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier16_Input2_10_0Output, mb_D_FF10_12MultiplierStage1Output);

    MB_D_FF_Float_10_12_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF10_12MultiplierStage1Output, mb_D_FF10_12MultiplierStage2Output);

    MB_D_FF_Float_Multiplier15_11_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier10_Output_12, mb_D_FFMultiplier15_11_0Output);

    MB_D_FF_Float_11_13_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier15_11_0Output, mb_D_FF11_13MultiplierStage1Output);

    MB_D_FF_Float_11_13_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF11_13MultiplierStage1Output, mb_D_FF11_13MultiplierStage2Output);

    Multiplier_Float_11: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF11_13MultiplierStage2Output, flopocoMultiplier11WeightInput, Multiplier11_Output_13);

    MBRightSHR_Float_11_13: entity work.MBRightSHR(rtl)
    GENERIC MAP (82, NumberOfBits)
    PORT MAP (clk, rst, Multiplier11Weight, mbRightSHR11_13Output);

    MB_D_FF_Float_11_13_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR11_13Output, Multiplier11WeightOutput);

    InputIEEE_Float_11_13: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier11WeightOutput, flopocoMultiplier11WeightOutput);

    MB_D_FF_Float_11_13_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier11WeightOutput, flopocoMultiplier11WeightInput);

    MBRightSHR_Float_12_Input114: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits)
    PORT MAP (clk, rst, Multiplier12Weight, mbRightSHR12_Input1_14Output);

    MB_D_FF_Float_12_14_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR12_Input1_14Output, Multiplier12WeightOutput);

    InputIEEE_Float_12_14: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier12WeightOutput, flopocoMultiplier12WeightOutput);

    MB_D_FF_Float_12_14_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier12WeightOutput, flopocoMultiplier12WeightInput);

    Multiplier_Float_12: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier12WeightInput, mb_D_FF12_14MultiplierStage2Output, Multiplier12_Output_14);

    MBRightSHR_Float_12_Input2_14: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR12_Input2_14Input, mbRightSHR12_Input2_14Output);

    MB_D_FF_Float_12_14_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR12_Input2_14Output, mb_D_FF12_14MultiplierStage1Output);

    MB_D_FF_Float_12_14_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF12_14MultiplierStage1Output, mb_D_FF12_14MultiplierStage2Output);

    MBRightSHR_Float_13_Input115: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits)
    PORT MAP (clk, rst, Multiplier13Weight, mbRightSHR13_Input1_15Output);

    MB_D_FF_Float_13_15_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR13_Input1_15Output, Multiplier13WeightOutput);

    InputIEEE_Float_13_15: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier13WeightOutput, flopocoMultiplier13WeightOutput);

    MB_D_FF_Float_13_15_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier13WeightOutput, flopocoMultiplier13WeightInput);

    Multiplier_Float_13: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier13WeightInput, mb_D_FF13_15MultiplierStage2Output, Multiplier13_Output_15);

    MBRightSHR_Float_13_Input2_15: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR13_Input2_15Input, mbRightSHR13_Input2_15Output);

    MB_D_FF_Float_13_15_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR13_Input2_15Output, mb_D_FF13_15MultiplierStage1Output);

    MB_D_FF_Float_13_15_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF13_15MultiplierStage1Output, mb_D_FF13_15MultiplierStage2Output);

    MB_D_FF_Float_Adder18_Input1_2_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier13_Output_15, mb_D_FFAdder18_Input1_2_0Output);

    MB_D_FF_Float_2_16_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder18_Input1_2_0Output, mb_D_FF2_16AugendStage1Output);

    MB_D_FF_Float_2_16_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF2_16AugendStage1Output, mb_D_FF2_16AugendStage2Output);

    Adder_Float_2: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF2_16AugendStage2Output, mb_D_FF2_16AddendStage2Output, Adder2_Output_16);

    MB_D_FF_Float_Adder18_Input2_2_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier12_Output_14, mb_D_FFAdder18_Input2_2_0Output);

    MB_D_FF_Float_2_16_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder18_Input2_2_0Output, mb_D_FF2_16AddendStage1Output);

    MB_D_FF_Float_2_16_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF2_16AddendStage1Output, mb_D_FF2_16AddendStage2Output);

    MB_D_FF_Float_Multiplier17_14_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder2_Output_16, mb_D_FFMultiplier17_14_0Output);

    MB_D_FF_Float_14_17_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier17_14_0Output, mb_D_FF14_17MultiplierStage1Output);

    MB_D_FF_Float_14_17_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF14_17MultiplierStage1Output, mb_D_FF14_17MultiplierStage2Output);

    Multiplier_Float_14: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF14_17MultiplierStage2Output, mb_D_FF14_17MultiplicandStage2Output, Multiplier14_Output_17);

    MBRightSHR_Float_14_17: entity work.MBRightSHR(rtl)
    GENERIC MAP (50, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR14_17Input, mbRightSHR14_17Output);

    MB_D_FF_Float_14_17_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR14_17Output, mb_D_FF14_17MultiplicandStage1Output);

    MB_D_FF_Float_14_17_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF14_17MultiplicandStage1Output, mb_D_FF14_17MultiplicandStage2Output);

    MB_D_FF_Float_Multiplier19_16_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier4_Output_5, mb_D_FFMultiplier19_16_0Output);

    MB_D_FF_Float_16_19_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier19_16_0Output, mb_D_FF16_19MultiplierStage1Output);

    MB_D_FF_Float_16_19_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF16_19MultiplierStage1Output, mb_D_FF16_19MultiplierStage2Output);

    Multiplier_Float_16: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF16_19MultiplierStage2Output, flopocoMultiplier16WeightInput, Multiplier16_Output_19);

    MBRightSHR_Float_16_19: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits)
    PORT MAP (clk, rst, Multiplier16Weight, mbRightSHR16_19Output);

    MB_D_FF_Float_16_19_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR16_19Output, Multiplier16WeightOutput);

    InputIEEE_Float_16_19: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier16WeightOutput, flopocoMultiplier16WeightOutput);

    MB_D_FF_Float_16_19_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier16WeightOutput, flopocoMultiplier16WeightInput);

    MB_D_FF_Float_Multiplier18_17_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier16_Output_19, mb_D_FFMultiplier18_17_0Output);

    MB_D_FF_Float_17_20_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier18_17_0Output, mb_D_FF17_20MultiplierStage1Output);

    MB_D_FF_Float_17_20_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF17_20MultiplierStage1Output, mb_D_FF17_20MultiplierStage2Output);

    Multiplier_Float_17: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF17_20MultiplierStage2Output, flopocoMultiplier17WeightInput, Multiplier17_Output_20);

    MBRightSHR_Float_17_20: entity work.MBRightSHR(rtl)
    GENERIC MAP (43, NumberOfBits)
    PORT MAP (clk, rst, Multiplier17Weight, mbRightSHR17_20Output);

    MB_D_FF_Float_17_20_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR17_20Output, Multiplier17WeightOutput);

    InputIEEE_Float_17_20: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier17WeightOutput, flopocoMultiplier17WeightOutput);

    MB_D_FF_Float_17_20_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier17WeightOutput, flopocoMultiplier17WeightInput);

    MB_D_FF_Float_Multiplier19_19_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier7_Output_8, mb_D_FFMultiplier19_19_0Output);

    MB_D_FF_Float_19_22_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier19_19_0Output, mb_D_FF19_22MultiplierStage1Output);

    MB_D_FF_Float_19_22_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF19_22MultiplierStage1Output, mb_D_FF19_22MultiplierStage2Output);

    Multiplier_Float_19: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF19_22MultiplierStage2Output, flopocoMultiplier19WeightInput, Multiplier19_Output_22);

    MBRightSHR_Float_19_22: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits)
    PORT MAP (clk, rst, Multiplier19Weight, mbRightSHR19_22Output);

    MB_D_FF_Float_19_22_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR19_22Output, Multiplier19WeightOutput);

    InputIEEE_Float_19_22: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier19WeightOutput, flopocoMultiplier19WeightOutput);

    MB_D_FF_Float_19_22_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier19WeightOutput, flopocoMultiplier19WeightInput);

    MB_D_FF_Float_Multiplier18_20_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier19_Output_22, mb_D_FFMultiplier18_20_0Output);

    MB_D_FF_Float_20_23_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier18_20_0Output, mb_D_FF20_23MultiplierStage1Output);

    MB_D_FF_Float_20_23_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF20_23MultiplierStage1Output, mb_D_FF20_23MultiplierStage2Output);

    Multiplier_Float_20: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF20_23MultiplierStage2Output, flopocoMultiplier20WeightInput, Multiplier20_Output_23);

    MBRightSHR_Float_20_23: entity work.MBRightSHR(rtl)
    GENERIC MAP (43, NumberOfBits)
    PORT MAP (clk, rst, Multiplier20Weight, mbRightSHR20_23Output);

    MB_D_FF_Float_20_23_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR20_23Output, Multiplier20WeightOutput);

    InputIEEE_Float_20_23: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier20WeightOutput, flopocoMultiplier20WeightOutput);

    MB_D_FF_Float_20_23_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier20WeightOutput, flopocoMultiplier20WeightInput);

    MB_D_FF_Float_Adder17_Input1_3_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier20_Output_23, mb_D_FFAdder17_Input1_3_0Output);

    MB_D_FF_Float_3_24_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder17_Input1_3_0Output, mb_D_FF3_24AugendStage1Output);

    MB_D_FF_Float_3_24_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF3_24AugendStage1Output, mb_D_FF3_24AugendStage2Output);

    Adder_Float_3: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF3_24AugendStage2Output, mb_D_FF3_24AddendStage2Output, Adder3_Output_24);

    MB_D_FF_Float_Adder17_Input2_3_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier17_Output_20, mb_D_FFAdder17_Input2_3_0Output);

    MB_D_FF_Float_3_24_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder17_Input2_3_0Output, mb_D_FF3_24AddendStage1Output);

    MB_D_FF_Float_3_24_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF3_24AddendStage1Output, mb_D_FF3_24AddendStage2Output);

    MB_D_FF_Float_Multiplier16_Input1_21_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder3_Output_24, mb_D_FFMultiplier16_Input1_21_0Output);

    MB_D_FF_Float_21_25_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier16_Input1_21_0Output, mb_D_FF21_25MultiplicandStage1Output);

    MB_D_FF_Float_21_25_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF21_25MultiplicandStage1Output, mb_D_FF21_25MultiplicandStage2Output);

    Multiplier_Float_21: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF21_25MultiplicandStage2Output, mb_D_FF21_25MultiplierStage2Output, Multiplier21_Output_25);

    MB_D_FF_Float_Multiplier16_Input2_21_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier14_Output_17, mb_D_FFMultiplier16_Input2_21_0Output);

    MB_D_FF_Float_21_25_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier16_Input2_21_0Output, mb_D_FF21_25MultiplierStage1Output);

    MB_D_FF_Float_21_25_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF21_25MultiplierStage1Output, mb_D_FF21_25MultiplierStage2Output);

    MB_D_FF_Float_Multiplier15_22_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier21_Output_25, mb_D_FFMultiplier15_22_0Output);

    MB_D_FF_Float_22_26_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier15_22_0Output, mb_D_FF22_26MultiplierStage1Output);

    MB_D_FF_Float_22_26_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF22_26MultiplierStage1Output, mb_D_FF22_26MultiplierStage2Output);

    Multiplier_Float_22: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF22_26MultiplierStage2Output, flopocoMultiplier22WeightInput, Multiplier22_Output_26);

    MBRightSHR_Float_22_26: entity work.MBRightSHR(rtl)
    GENERIC MAP (82, NumberOfBits)
    PORT MAP (clk, rst, Multiplier22Weight, mbRightSHR22_26Output);

    MB_D_FF_Float_22_26_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR22_26Output, Multiplier22WeightOutput);

    InputIEEE_Float_22_26: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier22WeightOutput, flopocoMultiplier22WeightOutput);

    MB_D_FF_Float_22_26_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier22WeightOutput, flopocoMultiplier22WeightInput);

    MB_D_FF_Float_Adder14_Input1_4_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier22_Output_26, mb_D_FFAdder14_Input1_4_0Output);

    MB_D_FF_Float_4_27_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder14_Input1_4_0Output, mb_D_FF4_27AugendStage1Output);

    MB_D_FF_Float_4_27_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF4_27AugendStage1Output, mb_D_FF4_27AugendStage2Output);

    Adder_Float_4: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF4_27AugendStage2Output, mb_D_FF4_27AddendStage2Output, Adder4_Output_27);

    MB_D_FF_Float_Adder14_Input2_4_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier11_Output_13, mb_D_FFAdder14_Input2_4_0Output);

    MB_D_FF_Float_4_27_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder14_Input2_4_0Output, mb_D_FF4_27AddendStage1Output);

    MB_D_FF_Float_4_27_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF4_27AddendStage1Output, mb_D_FF4_27AddendStage2Output);

    MB_D_FF_Float_Multiplier13_Input1_23_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder4_Output_27, mb_D_FFMultiplier13_Input1_23_0Output);

    MB_D_FF_Float_23_28_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier13_Input1_23_0Output, mb_D_FF23_28MultiplicandStage1Output);

    MB_D_FF_Float_23_28_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF23_28MultiplicandStage1Output, mb_D_FF23_28MultiplicandStage2Output);

    Multiplier_Float_23: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF23_28MultiplicandStage2Output, mb_D_FF23_28MultiplierStage2Output, Multiplier23_Output_28);

    MB_D_FF_Float_Multiplier13_Input2_23_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier0_Output_0, mb_D_FFMultiplier13_Input2_23_0Output);

    MB_D_FF_Float_23_28_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier13_Input2_23_0Output, mb_D_FF23_28MultiplierStage1Output);

    MB_D_FF_Float_23_28_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF23_28MultiplierStage1Output, mb_D_FF23_28MultiplierStage2Output);

    MB_D_FF_Float_Multiplier12_24_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier23_Output_28, mb_D_FFMultiplier12_24_0Output);

    MB_D_FF_Float_24_29_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier12_24_0Output, mb_D_FF24_29MultiplierStage1Output);

    MB_D_FF_Float_24_29_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF24_29MultiplierStage1Output, mb_D_FF24_29MultiplierStage2Output);

    Multiplier_Float_24: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF24_29MultiplierStage2Output, flopocoMultiplier24WeightInput, Multiplier24_Output_29);

    MBRightSHR_Float_24_29: entity work.MBRightSHR(rtl)
    GENERIC MAP (121, NumberOfBits)
    PORT MAP (clk, rst, Multiplier24Weight, mbRightSHR24_29Output);

    MB_D_FF_Float_24_29_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR24_29Output, Multiplier24WeightOutput);

    InputIEEE_Float_24_29: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier24WeightOutput, flopocoMultiplier24WeightOutput);

    MB_D_FF_Float_24_29_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier24WeightOutput, flopocoMultiplier24WeightInput);

    MBRightSHR_Float_25_Input130: entity work.MBRightSHR(rtl)
    GENERIC MAP (89, NumberOfBits)
    PORT MAP (clk, rst, Multiplier25Weight, mbRightSHR25_Input1_30Output);

    MB_D_FF_Float_25_30_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR25_Input1_30Output, Multiplier25WeightOutput);

    InputIEEE_Float_25_30: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier25WeightOutput, flopocoMultiplier25WeightOutput);

    MB_D_FF_Float_25_30_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier25WeightOutput, flopocoMultiplier25WeightInput);

    Multiplier_Float_25: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier25WeightInput, mb_D_FF25_30MultiplierStage2Output, Multiplier25_Output_30);

    MBRightSHR_Float_25_Input2_30: entity work.MBRightSHR(rtl)
    GENERIC MAP (89, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR25_Input2_30Input, mbRightSHR25_Input2_30Output);

    MB_D_FF_Float_25_30_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR25_Input2_30Output, mb_D_FF25_30MultiplierStage1Output);

    MB_D_FF_Float_25_30_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF25_30MultiplierStage1Output, mb_D_FF25_30MultiplierStage2Output);

    MBRightSHR_Float_26_Input131: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits)
    PORT MAP (clk, rst, Multiplier26Weight, mbRightSHR26_Input1_31Output);

    MB_D_FF_Float_26_31_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR26_Input1_31Output, Multiplier26WeightOutput);

    InputIEEE_Float_26_31: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier26WeightOutput, flopocoMultiplier26WeightOutput);

    MB_D_FF_Float_26_31_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier26WeightOutput, flopocoMultiplier26WeightInput);

    Multiplier_Float_26: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier26WeightInput, mb_D_FF26_31MultiplierStage2Output, Multiplier26_Output_31);

    MBRightSHR_Float_26_Input2_31: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR26_Input2_31Input, mbRightSHR26_Input2_31Output);

    MB_D_FF_Float_26_31_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR26_Input2_31Output, mb_D_FF26_31MultiplierStage1Output);

    MB_D_FF_Float_26_31_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF26_31MultiplierStage1Output, mb_D_FF26_31MultiplierStage2Output);

    MBRightSHR_Float_27_Input132: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits)
    PORT MAP (clk, rst, Multiplier27Weight, mbRightSHR27_Input1_32Output);

    MB_D_FF_Float_27_32_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR27_Input1_32Output, Multiplier27WeightOutput);

    InputIEEE_Float_27_32: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier27WeightOutput, flopocoMultiplier27WeightOutput);

    MB_D_FF_Float_27_32_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier27WeightOutput, flopocoMultiplier27WeightInput);

    Multiplier_Float_27: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier27WeightInput, mb_D_FF27_32MultiplierStage2Output, Multiplier27_Output_32);

    MBRightSHR_Float_27_Input2_32: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR27_Input2_32Input, mbRightSHR27_Input2_32Output);

    MB_D_FF_Float_27_32_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR27_Input2_32Output, mb_D_FF27_32MultiplierStage1Output);

    MB_D_FF_Float_27_32_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF27_32MultiplierStage1Output, mb_D_FF27_32MultiplierStage2Output);

    MB_D_FF_Float_Adder18_Input1_5_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier27_Output_32, mb_D_FFAdder18_Input1_5_0Output);

    MB_D_FF_Float_5_33_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder18_Input1_5_0Output, mb_D_FF5_33AugendStage1Output);

    MB_D_FF_Float_5_33_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF5_33AugendStage1Output, mb_D_FF5_33AugendStage2Output);

    Adder_Float_5: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF5_33AugendStage2Output, mb_D_FF5_33AddendStage2Output, Adder5_Output_33);

    MB_D_FF_Float_Adder18_Input2_5_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier26_Output_31, mb_D_FFAdder18_Input2_5_0Output);

    MB_D_FF_Float_5_33_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder18_Input2_5_0Output, mb_D_FF5_33AddendStage1Output);

    MB_D_FF_Float_5_33_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF5_33AddendStage1Output, mb_D_FF5_33AddendStage2Output);

    MB_D_FF_Float_Multiplier17_28_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder5_Output_33, mb_D_FFMultiplier17_28_0Output);

    MB_D_FF_Float_28_34_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier17_28_0Output, mb_D_FF28_34MultiplierStage1Output);

    MB_D_FF_Float_28_34_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF28_34MultiplierStage1Output, mb_D_FF28_34MultiplierStage2Output);

    Multiplier_Float_28: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF28_34MultiplierStage2Output, mb_D_FF28_34MultiplicandStage2Output, Multiplier28_Output_34);

    MBRightSHR_Float_28_34: entity work.MBRightSHR(rtl)
    GENERIC MAP (50, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR28_34Input, mbRightSHR28_34Output);

    MB_D_FF_Float_28_34_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR28_34Output, mb_D_FF28_34MultiplicandStage1Output);

    MB_D_FF_Float_28_34_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF28_34MultiplicandStage1Output, mb_D_FF28_34MultiplicandStage2Output);

    MBRightSHR_Float_29_Input135: entity work.MBRightSHR(rtl)
    GENERIC MAP (11, NumberOfBits)
    PORT MAP (clk, rst, Multiplier29Weight, mbRightSHR29_Input1_35Output);

    MB_D_FF_Float_29_35_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR29_Input1_35Output, Multiplier29WeightOutput);

    InputIEEE_Float_29_35: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier29WeightOutput, flopocoMultiplier29WeightOutput);

    MB_D_FF_Float_29_35_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier29WeightOutput, flopocoMultiplier29WeightInput);

    Multiplier_Float_29: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier29WeightInput, mb_D_FF29_35MultiplierStage2Output, Multiplier29_Output_35);

    MBRightSHR_Float_29_Input2_35: entity work.MBRightSHR(rtl)
    GENERIC MAP (11, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR29_Input2_35Input, mbRightSHR29_Input2_35Output);

    MB_D_FF_Float_29_35_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR29_Input2_35Output, mb_D_FF29_35MultiplierStage1Output);

    MB_D_FF_Float_29_35_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF29_35MultiplierStage1Output, mb_D_FF29_35MultiplierStage2Output);

    MB_D_FF_Float_Multiplier19_30_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier29_Output_35, mb_D_FFMultiplier19_30_0Output);

    MB_D_FF_Float_30_36_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier19_30_0Output, mb_D_FF30_36MultiplierStage1Output);

    MB_D_FF_Float_30_36_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF30_36MultiplierStage1Output, mb_D_FF30_36MultiplierStage2Output);

    Multiplier_Float_30: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF30_36MultiplierStage2Output, flopocoMultiplier30WeightInput, Multiplier30_Output_36);

    MBRightSHR_Float_30_36: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits)
    PORT MAP (clk, rst, Multiplier30Weight, mbRightSHR30_36Output);

    MB_D_FF_Float_30_36_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR30_36Output, Multiplier30WeightOutput);

    InputIEEE_Float_30_36: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier30WeightOutput, flopocoMultiplier30WeightOutput);

    MB_D_FF_Float_30_36_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier30WeightOutput, flopocoMultiplier30WeightInput);

    MB_D_FF_Float_Multiplier18_31_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier30_Output_36, mb_D_FFMultiplier18_31_0Output);

    MB_D_FF_Float_31_37_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier18_31_0Output, mb_D_FF31_37MultiplierStage1Output);

    MB_D_FF_Float_31_37_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF31_37MultiplierStage1Output, mb_D_FF31_37MultiplierStage2Output);

    Multiplier_Float_31: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF31_37MultiplierStage2Output, flopocoMultiplier31WeightInput, Multiplier31_Output_37);

    MBRightSHR_Float_31_37: entity work.MBRightSHR(rtl)
    GENERIC MAP (43, NumberOfBits)
    PORT MAP (clk, rst, Multiplier31Weight, mbRightSHR31_37Output);

    MB_D_FF_Float_31_37_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR31_37Output, Multiplier31WeightOutput);

    InputIEEE_Float_31_37: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier31WeightOutput, flopocoMultiplier31WeightOutput);

    MB_D_FF_Float_31_37_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier31WeightOutput, flopocoMultiplier31WeightInput);

    MBRightSHR_Float_32_Input138: entity work.MBRightSHR(rtl)
    GENERIC MAP (11, NumberOfBits)
    PORT MAP (clk, rst, Multiplier32Weight, mbRightSHR32_Input1_38Output);

    MB_D_FF_Float_32_38_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR32_Input1_38Output, Multiplier32WeightOutput);

    InputIEEE_Float_32_38: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier32WeightOutput, flopocoMultiplier32WeightOutput);

    MB_D_FF_Float_32_38_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier32WeightOutput, flopocoMultiplier32WeightInput);

    Multiplier_Float_32: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier32WeightInput, mb_D_FF32_38MultiplierStage2Output, Multiplier32_Output_38);

    MBRightSHR_Float_32_Input2_38: entity work.MBRightSHR(rtl)
    GENERIC MAP (11, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR32_Input2_38Input, mbRightSHR32_Input2_38Output);

    MB_D_FF_Float_32_38_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR32_Input2_38Output, mb_D_FF32_38MultiplierStage1Output);

    MB_D_FF_Float_32_38_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF32_38MultiplierStage1Output, mb_D_FF32_38MultiplierStage2Output);

    MB_D_FF_Float_Multiplier19_33_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier32_Output_38, mb_D_FFMultiplier19_33_0Output);

    MB_D_FF_Float_33_39_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier19_33_0Output, mb_D_FF33_39MultiplierStage1Output);

    MB_D_FF_Float_33_39_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF33_39MultiplierStage1Output, mb_D_FF33_39MultiplierStage2Output);

    Multiplier_Float_33: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF33_39MultiplierStage2Output, flopocoMultiplier33WeightInput, Multiplier33_Output_39);

    MBRightSHR_Float_33_39: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits)
    PORT MAP (clk, rst, Multiplier33Weight, mbRightSHR33_39Output);

    MB_D_FF_Float_33_39_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR33_39Output, Multiplier33WeightOutput);

    InputIEEE_Float_33_39: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier33WeightOutput, flopocoMultiplier33WeightOutput);

    MB_D_FF_Float_33_39_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier33WeightOutput, flopocoMultiplier33WeightInput);

    MB_D_FF_Float_Multiplier18_34_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier33_Output_39, mb_D_FFMultiplier18_34_0Output);

    MB_D_FF_Float_34_40_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier18_34_0Output, mb_D_FF34_40MultiplierStage1Output);

    MB_D_FF_Float_34_40_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF34_40MultiplierStage1Output, mb_D_FF34_40MultiplierStage2Output);

    Multiplier_Float_34: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF34_40MultiplierStage2Output, flopocoMultiplier34WeightInput, Multiplier34_Output_40);

    MBRightSHR_Float_34_40: entity work.MBRightSHR(rtl)
    GENERIC MAP (43, NumberOfBits)
    PORT MAP (clk, rst, Multiplier34Weight, mbRightSHR34_40Output);

    MB_D_FF_Float_34_40_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR34_40Output, Multiplier34WeightOutput);

    InputIEEE_Float_34_40: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier34WeightOutput, flopocoMultiplier34WeightOutput);

    MB_D_FF_Float_34_40_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier34WeightOutput, flopocoMultiplier34WeightInput);

    MB_D_FF_Float_Adder17_Input1_6_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier34_Output_40, mb_D_FFAdder17_Input1_6_0Output);

    MB_D_FF_Float_6_41_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder17_Input1_6_0Output, mb_D_FF6_41AugendStage1Output);

    MB_D_FF_Float_6_41_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF6_41AugendStage1Output, mb_D_FF6_41AugendStage2Output);

    Adder_Float_6: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF6_41AugendStage2Output, mb_D_FF6_41AddendStage2Output, Adder6_Output_41);

    MB_D_FF_Float_Adder17_Input2_6_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier31_Output_37, mb_D_FFAdder17_Input2_6_0Output);

    MB_D_FF_Float_6_41_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder17_Input2_6_0Output, mb_D_FF6_41AddendStage1Output);

    MB_D_FF_Float_6_41_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF6_41AddendStage1Output, mb_D_FF6_41AddendStage2Output);

    MB_D_FF_Float_Multiplier16_Input1_35_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder6_Output_41, mb_D_FFMultiplier16_Input1_35_0Output);

    MB_D_FF_Float_35_42_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier16_Input1_35_0Output, mb_D_FF35_42MultiplicandStage1Output);

    MB_D_FF_Float_35_42_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF35_42MultiplicandStage1Output, mb_D_FF35_42MultiplicandStage2Output);

    Multiplier_Float_35: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF35_42MultiplicandStage2Output, mb_D_FF35_42MultiplierStage2Output, Multiplier35_Output_42);

    MB_D_FF_Float_Multiplier16_Input2_35_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier28_Output_34, mb_D_FFMultiplier16_Input2_35_0Output);

    MB_D_FF_Float_35_42_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier16_Input2_35_0Output, mb_D_FF35_42MultiplierStage1Output);

    MB_D_FF_Float_35_42_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF35_42MultiplierStage1Output, mb_D_FF35_42MultiplierStage2Output);

    MB_D_FF_Float_Multiplier15_36_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier35_Output_42, mb_D_FFMultiplier15_36_0Output);

    MB_D_FF_Float_36_43_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier15_36_0Output, mb_D_FF36_43MultiplierStage1Output);

    MB_D_FF_Float_36_43_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF36_43MultiplierStage1Output, mb_D_FF36_43MultiplierStage2Output);

    Multiplier_Float_36: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF36_43MultiplierStage2Output, flopocoMultiplier36WeightInput, Multiplier36_Output_43);

    MBRightSHR_Float_36_43: entity work.MBRightSHR(rtl)
    GENERIC MAP (82, NumberOfBits)
    PORT MAP (clk, rst, Multiplier36Weight, mbRightSHR36_43Output);

    MB_D_FF_Float_36_43_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR36_43Output, Multiplier36WeightOutput);

    InputIEEE_Float_36_43: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier36WeightOutput, flopocoMultiplier36WeightOutput);

    MB_D_FF_Float_36_43_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier36WeightOutput, flopocoMultiplier36WeightInput);

    MBRightSHR_Float_37_Input144: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits)
    PORT MAP (clk, rst, Multiplier37Weight, mbRightSHR37_Input1_44Output);

    MB_D_FF_Float_37_44_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR37_Input1_44Output, Multiplier37WeightOutput);

    InputIEEE_Float_37_44: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier37WeightOutput, flopocoMultiplier37WeightOutput);

    MB_D_FF_Float_37_44_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier37WeightOutput, flopocoMultiplier37WeightInput);

    Multiplier_Float_37: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier37WeightInput, mb_D_FF37_44MultiplierStage2Output, Multiplier37_Output_44);

    MBRightSHR_Float_37_Input2_44: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR37_Input2_44Input, mbRightSHR37_Input2_44Output);

    MB_D_FF_Float_37_44_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR37_Input2_44Output, mb_D_FF37_44MultiplierStage1Output);

    MB_D_FF_Float_37_44_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF37_44MultiplierStage1Output, mb_D_FF37_44MultiplierStage2Output);

    MBRightSHR_Float_38_Input145: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits)
    PORT MAP (clk, rst, Multiplier38Weight, mbRightSHR38_Input1_45Output);

    MB_D_FF_Float_38_45_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR38_Input1_45Output, Multiplier38WeightOutput);

    InputIEEE_Float_38_45: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier38WeightOutput, flopocoMultiplier38WeightOutput);

    MB_D_FF_Float_38_45_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier38WeightOutput, flopocoMultiplier38WeightInput);

    Multiplier_Float_38: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier38WeightInput, mb_D_FF38_45MultiplierStage2Output, Multiplier38_Output_45);

    MBRightSHR_Float_38_Input2_45: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR38_Input2_45Input, mbRightSHR38_Input2_45Output);

    MB_D_FF_Float_38_45_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR38_Input2_45Output, mb_D_FF38_45MultiplierStage1Output);

    MB_D_FF_Float_38_45_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF38_45MultiplierStage1Output, mb_D_FF38_45MultiplierStage2Output);

    MB_D_FF_Float_Adder18_Input1_7_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier38_Output_45, mb_D_FFAdder18_Input1_7_0Output);

    MB_D_FF_Float_7_46_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder18_Input1_7_0Output, mb_D_FF7_46AugendStage1Output);

    MB_D_FF_Float_7_46_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF7_46AugendStage1Output, mb_D_FF7_46AugendStage2Output);

    Adder_Float_7: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF7_46AugendStage2Output, mb_D_FF7_46AddendStage2Output, Adder7_Output_46);

    MB_D_FF_Float_Adder18_Input2_7_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier37_Output_44, mb_D_FFAdder18_Input2_7_0Output);

    MB_D_FF_Float_7_46_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder18_Input2_7_0Output, mb_D_FF7_46AddendStage1Output);

    MB_D_FF_Float_7_46_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF7_46AddendStage1Output, mb_D_FF7_46AddendStage2Output);

    MB_D_FF_Float_Multiplier17_39_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder7_Output_46, mb_D_FFMultiplier17_39_0Output);

    MB_D_FF_Float_39_47_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier17_39_0Output, mb_D_FF39_47MultiplierStage1Output);

    MB_D_FF_Float_39_47_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF39_47MultiplierStage1Output, mb_D_FF39_47MultiplierStage2Output);

    Multiplier_Float_39: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF39_47MultiplierStage2Output, mb_D_FF39_47MultiplicandStage2Output, Multiplier39_Output_47);

    MBRightSHR_Float_39_47: entity work.MBRightSHR(rtl)
    GENERIC MAP (50, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR39_47Input, mbRightSHR39_47Output);

    MB_D_FF_Float_39_47_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR39_47Output, mb_D_FF39_47MultiplicandStage1Output);

    MB_D_FF_Float_39_47_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF39_47MultiplicandStage1Output, mb_D_FF39_47MultiplicandStage2Output);

    MB_D_FF_Float_Multiplier19_41_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier29_Output_35, mb_D_FFMultiplier19_41_0Output);

    MB_D_FF_Float_41_49_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier19_41_0Output, mb_D_FF41_49MultiplierStage1Output);

    MB_D_FF_Float_41_49_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF41_49MultiplierStage1Output, mb_D_FF41_49MultiplierStage2Output);

    Multiplier_Float_41: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF41_49MultiplierStage2Output, flopocoMultiplier41WeightInput, Multiplier41_Output_49);

    MBRightSHR_Float_41_49: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits)
    PORT MAP (clk, rst, Multiplier41Weight, mbRightSHR41_49Output);

    MB_D_FF_Float_41_49_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR41_49Output, Multiplier41WeightOutput);

    InputIEEE_Float_41_49: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier41WeightOutput, flopocoMultiplier41WeightOutput);

    MB_D_FF_Float_41_49_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier41WeightOutput, flopocoMultiplier41WeightInput);

    MB_D_FF_Float_Multiplier18_42_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier41_Output_49, mb_D_FFMultiplier18_42_0Output);

    MB_D_FF_Float_42_50_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier18_42_0Output, mb_D_FF42_50MultiplierStage1Output);

    MB_D_FF_Float_42_50_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF42_50MultiplierStage1Output, mb_D_FF42_50MultiplierStage2Output);

    Multiplier_Float_42: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF42_50MultiplierStage2Output, flopocoMultiplier42WeightInput, Multiplier42_Output_50);

    MBRightSHR_Float_42_50: entity work.MBRightSHR(rtl)
    GENERIC MAP (43, NumberOfBits)
    PORT MAP (clk, rst, Multiplier42Weight, mbRightSHR42_50Output);

    MB_D_FF_Float_42_50_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR42_50Output, Multiplier42WeightOutput);

    InputIEEE_Float_42_50: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier42WeightOutput, flopocoMultiplier42WeightOutput);

    MB_D_FF_Float_42_50_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier42WeightOutput, flopocoMultiplier42WeightInput);

    MB_D_FF_Float_Multiplier19_44_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier32_Output_38, mb_D_FFMultiplier19_44_0Output);

    MB_D_FF_Float_44_52_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier19_44_0Output, mb_D_FF44_52MultiplierStage1Output);

    MB_D_FF_Float_44_52_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF44_52MultiplierStage1Output, mb_D_FF44_52MultiplierStage2Output);

    Multiplier_Float_44: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF44_52MultiplierStage2Output, flopocoMultiplier44WeightInput, Multiplier44_Output_52);

    MBRightSHR_Float_44_52: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits)
    PORT MAP (clk, rst, Multiplier44Weight, mbRightSHR44_52Output);

    MB_D_FF_Float_44_52_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR44_52Output, Multiplier44WeightOutput);

    InputIEEE_Float_44_52: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier44WeightOutput, flopocoMultiplier44WeightOutput);

    MB_D_FF_Float_44_52_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier44WeightOutput, flopocoMultiplier44WeightInput);

    MB_D_FF_Float_Multiplier18_45_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier44_Output_52, mb_D_FFMultiplier18_45_0Output);

    MB_D_FF_Float_45_53_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier18_45_0Output, mb_D_FF45_53MultiplierStage1Output);

    MB_D_FF_Float_45_53_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF45_53MultiplierStage1Output, mb_D_FF45_53MultiplierStage2Output);

    Multiplier_Float_45: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF45_53MultiplierStage2Output, flopocoMultiplier45WeightInput, Multiplier45_Output_53);

    MBRightSHR_Float_45_53: entity work.MBRightSHR(rtl)
    GENERIC MAP (43, NumberOfBits)
    PORT MAP (clk, rst, Multiplier45Weight, mbRightSHR45_53Output);

    MB_D_FF_Float_45_53_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR45_53Output, Multiplier45WeightOutput);

    InputIEEE_Float_45_53: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier45WeightOutput, flopocoMultiplier45WeightOutput);

    MB_D_FF_Float_45_53_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier45WeightOutput, flopocoMultiplier45WeightInput);

    MB_D_FF_Float_Adder17_Input1_8_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier45_Output_53, mb_D_FFAdder17_Input1_8_0Output);

    MB_D_FF_Float_8_54_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder17_Input1_8_0Output, mb_D_FF8_54AugendStage1Output);

    MB_D_FF_Float_8_54_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF8_54AugendStage1Output, mb_D_FF8_54AugendStage2Output);

    Adder_Float_8: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF8_54AugendStage2Output, mb_D_FF8_54AddendStage2Output, Adder8_Output_54);

    MB_D_FF_Float_Adder17_Input2_8_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier42_Output_50, mb_D_FFAdder17_Input2_8_0Output);

    MB_D_FF_Float_8_54_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder17_Input2_8_0Output, mb_D_FF8_54AddendStage1Output);

    MB_D_FF_Float_8_54_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF8_54AddendStage1Output, mb_D_FF8_54AddendStage2Output);

    MB_D_FF_Float_Multiplier16_Input1_46_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder8_Output_54, mb_D_FFMultiplier16_Input1_46_0Output);

    MB_D_FF_Float_46_55_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier16_Input1_46_0Output, mb_D_FF46_55MultiplicandStage1Output);

    MB_D_FF_Float_46_55_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF46_55MultiplicandStage1Output, mb_D_FF46_55MultiplicandStage2Output);

    Multiplier_Float_46: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF46_55MultiplicandStage2Output, mb_D_FF46_55MultiplierStage2Output, Multiplier46_Output_55);

    MB_D_FF_Float_Multiplier16_Input2_46_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier39_Output_47, mb_D_FFMultiplier16_Input2_46_0Output);

    MB_D_FF_Float_46_55_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier16_Input2_46_0Output, mb_D_FF46_55MultiplierStage1Output);

    MB_D_FF_Float_46_55_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF46_55MultiplierStage1Output, mb_D_FF46_55MultiplierStage2Output);

    MB_D_FF_Float_Multiplier15_47_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier46_Output_55, mb_D_FFMultiplier15_47_0Output);

    MB_D_FF_Float_47_56_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier15_47_0Output, mb_D_FF47_56MultiplierStage1Output);

    MB_D_FF_Float_47_56_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF47_56MultiplierStage1Output, mb_D_FF47_56MultiplierStage2Output);

    Multiplier_Float_47: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF47_56MultiplierStage2Output, flopocoMultiplier47WeightInput, Multiplier47_Output_56);

    MBRightSHR_Float_47_56: entity work.MBRightSHR(rtl)
    GENERIC MAP (82, NumberOfBits)
    PORT MAP (clk, rst, Multiplier47Weight, mbRightSHR47_56Output);

    MB_D_FF_Float_47_56_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR47_56Output, Multiplier47WeightOutput);

    InputIEEE_Float_47_56: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier47WeightOutput, flopocoMultiplier47WeightOutput);

    MB_D_FF_Float_47_56_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier47WeightOutput, flopocoMultiplier47WeightInput);

    MB_D_FF_Float_Adder14_Input1_9_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier47_Output_56, mb_D_FFAdder14_Input1_9_0Output);

    MB_D_FF_Float_9_57_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder14_Input1_9_0Output, mb_D_FF9_57AugendStage1Output);

    MB_D_FF_Float_9_57_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF9_57AugendStage1Output, mb_D_FF9_57AugendStage2Output);

    Adder_Float_9: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF9_57AugendStage2Output, mb_D_FF9_57AddendStage2Output, Adder9_Output_57);

    MB_D_FF_Float_Adder14_Input2_9_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier36_Output_43, mb_D_FFAdder14_Input2_9_0Output);

    MB_D_FF_Float_9_57_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder14_Input2_9_0Output, mb_D_FF9_57AddendStage1Output);

    MB_D_FF_Float_9_57_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF9_57AddendStage1Output, mb_D_FF9_57AddendStage2Output);

    MB_D_FF_Float_Multiplier13_Input1_48_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder9_Output_57, mb_D_FFMultiplier13_Input1_48_0Output);

    MB_D_FF_Float_48_58_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier13_Input1_48_0Output, mb_D_FF48_58MultiplicandStage1Output);

    MB_D_FF_Float_48_58_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF48_58MultiplicandStage1Output, mb_D_FF48_58MultiplicandStage2Output);

    Multiplier_Float_48: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF48_58MultiplicandStage2Output, mb_D_FF48_58MultiplierStage2Output, Multiplier48_Output_58);

    MB_D_FF_Float_Multiplier13_Input2_48_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier25_Output_30, mb_D_FFMultiplier13_Input2_48_0Output);

    MB_D_FF_Float_48_58_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier13_Input2_48_0Output, mb_D_FF48_58MultiplierStage1Output);

    MB_D_FF_Float_48_58_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF48_58MultiplierStage1Output, mb_D_FF48_58MultiplierStage2Output);

    MB_D_FF_Float_Multiplier12_49_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier48_Output_58, mb_D_FFMultiplier12_49_0Output);

    MB_D_FF_Float_49_59_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier12_49_0Output, mb_D_FF49_59MultiplierStage1Output);

    MB_D_FF_Float_49_59_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF49_59MultiplierStage1Output, mb_D_FF49_59MultiplierStage2Output);

    Multiplier_Float_49: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF49_59MultiplierStage2Output, flopocoMultiplier49WeightInput, Multiplier49_Output_59);

    MBRightSHR_Float_49_59: entity work.MBRightSHR(rtl)
    GENERIC MAP (121, NumberOfBits)
    PORT MAP (clk, rst, Multiplier49Weight, mbRightSHR49_59Output);

    MB_D_FF_Float_49_59_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR49_59Output, Multiplier49WeightOutput);

    InputIEEE_Float_49_59: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier49WeightOutput, flopocoMultiplier49WeightOutput);

    MB_D_FF_Float_49_59_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier49WeightOutput, flopocoMultiplier49WeightInput);

    MB_D_FF_Float_Adder11_Input1_10_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier49_Output_59, mb_D_FFAdder11_Input1_10_0Output);

    MB_D_FF_Float_10_60_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder11_Input1_10_0Output, mb_D_FF10_60AugendStage1Output);

    MB_D_FF_Float_10_60_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF10_60AugendStage1Output, mb_D_FF10_60AugendStage2Output);

    Adder_Float_10: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF10_60AugendStage2Output, mb_D_FF10_60AddendStage2Output, Adder10_Output_60);

    MB_D_FF_Float_Adder11_Input2_10_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier24_Output_29, mb_D_FFAdder11_Input2_10_0Output);

    MB_D_FF_Float_10_60_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder11_Input2_10_0Output, mb_D_FF10_60AddendStage1Output);

    MB_D_FF_Float_10_60_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF10_60AddendStage1Output, mb_D_FF10_60AddendStage2Output);

    MB_D_FF_Float_Multiplier10_50_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder10_Output_60, mb_D_FFMultiplier10_50_0Output);

    MB_D_FF_Float_50_61_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier10_50_0Output, mb_D_FF50_61MultiplierStage1Output);

    MB_D_FF_Float_50_61_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF50_61MultiplierStage1Output, mb_D_FF50_61MultiplierStage2Output);

    Multiplier_Float_50: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF50_61MultiplierStage2Output, mb_D_FF50_61MultiplicandStage2Output, Multiplier50_Output_61);

    MBRightSHR_Float_50_61: entity work.MBRightSHR(rtl)
    GENERIC MAP (135, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR50_61Input, mbRightSHR50_61Output);

    MB_D_FF_Float_50_61_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR50_61Output, mb_D_FF50_61MultiplicandStage1Output);

    MB_D_FF_Float_50_61_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF50_61MultiplicandStage1Output, mb_D_FF50_61MultiplicandStage2Output);

    MB_D_FF_Float_Multiplier9_51_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier50_Output_61, mb_D_FFMultiplier9_51_0Output);

    MB_D_FF_Float_51_62_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier9_51_0Output, mb_D_FF51_62MultiplierStage1Output);

    MB_D_FF_Float_51_62_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF51_62MultiplierStage1Output, mb_D_FF51_62MultiplierStage2Output);

    Multiplier_Float_51: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF51_62MultiplierStage2Output, flopocoMultiplier51WeightInput, Multiplier51_Output_62);

    MBRightSHR_Float_51_62: entity work.MBRightSHR(rtl)
    GENERIC MAP (160, NumberOfBits)
    PORT MAP (clk, rst, Multiplier51Weight, mbRightSHR51_62Output);

    MB_D_FF_Float_51_62_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR51_62Output, Multiplier51WeightOutput);

    InputIEEE_Float_51_62: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier51WeightOutput, flopocoMultiplier51WeightOutput);

    MB_D_FF_Float_51_62_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier51WeightOutput, flopocoMultiplier51WeightInput);

    MBRightSHR_Float_53_Input164: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits)
    PORT MAP (clk, rst, Multiplier53Weight, mbRightSHR53_Input1_64Output);

    MB_D_FF_Float_53_64_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR53_Input1_64Output, Multiplier53WeightOutput);

    InputIEEE_Float_53_64: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier53WeightOutput, flopocoMultiplier53WeightOutput);

    MB_D_FF_Float_53_64_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier53WeightOutput, flopocoMultiplier53WeightInput);

    Multiplier_Float_53: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier53WeightInput, mb_D_FF53_64MultiplierStage2Output, Multiplier53_Output_64);

    MBRightSHR_Float_53_Input2_64: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR53_Input2_64Input, mbRightSHR53_Input2_64Output);

    MB_D_FF_Float_53_64_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR53_Input2_64Output, mb_D_FF53_64MultiplierStage1Output);

    MB_D_FF_Float_53_64_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF53_64MultiplierStage1Output, mb_D_FF53_64MultiplierStage2Output);

    MBRightSHR_Float_54_Input165: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits)
    PORT MAP (clk, rst, Multiplier54Weight, mbRightSHR54_Input1_65Output);

    MB_D_FF_Float_54_65_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR54_Input1_65Output, Multiplier54WeightOutput);

    InputIEEE_Float_54_65: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier54WeightOutput, flopocoMultiplier54WeightOutput);

    MB_D_FF_Float_54_65_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier54WeightOutput, flopocoMultiplier54WeightInput);

    Multiplier_Float_54: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier54WeightInput, mb_D_FF54_65MultiplierStage2Output, Multiplier54_Output_65);

    MBRightSHR_Float_54_Input2_65: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR54_Input2_65Input, mbRightSHR54_Input2_65Output);

    MB_D_FF_Float_54_65_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR54_Input2_65Output, mb_D_FF54_65MultiplierStage1Output);

    MB_D_FF_Float_54_65_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF54_65MultiplierStage1Output, mb_D_FF54_65MultiplierStage2Output);

    MB_D_FF_Float_Adder18_Input1_11_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier54_Output_65, mb_D_FFAdder18_Input1_11_0Output);

    MB_D_FF_Float_11_66_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder18_Input1_11_0Output, mb_D_FF11_66AugendStage1Output);

    MB_D_FF_Float_11_66_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF11_66AugendStage1Output, mb_D_FF11_66AugendStage2Output);

    Adder_Float_11: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF11_66AugendStage2Output, mb_D_FF11_66AddendStage2Output, Adder11_Output_66);

    MB_D_FF_Float_Adder18_Input2_11_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier53_Output_64, mb_D_FFAdder18_Input2_11_0Output);

    MB_D_FF_Float_11_66_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder18_Input2_11_0Output, mb_D_FF11_66AddendStage1Output);

    MB_D_FF_Float_11_66_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF11_66AddendStage1Output, mb_D_FF11_66AddendStage2Output);

    MB_D_FF_Float_Multiplier17_55_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder11_Output_66, mb_D_FFMultiplier17_55_0Output);

    MB_D_FF_Float_55_67_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier17_55_0Output, mb_D_FF55_67MultiplierStage1Output);

    MB_D_FF_Float_55_67_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF55_67MultiplierStage1Output, mb_D_FF55_67MultiplierStage2Output);

    Multiplier_Float_55: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF55_67MultiplierStage2Output, mb_D_FF55_67MultiplicandStage2Output, Multiplier55_Output_67);

    MBRightSHR_Float_55_67: entity work.MBRightSHR(rtl)
    GENERIC MAP (50, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR55_67Input, mbRightSHR55_67Output);

    MB_D_FF_Float_55_67_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR55_67Output, mb_D_FF55_67MultiplicandStage1Output);

    MB_D_FF_Float_55_67_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF55_67MultiplicandStage1Output, mb_D_FF55_67MultiplicandStage2Output);

    MB_D_FF_Float_Multiplier18_58_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier5_Output_6, mb_D_FFMultiplier18_58_0Output);

    MB_D_FF_Float_58_70_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier18_58_0Output, mb_D_FF58_70MultiplierStage1Output);

    MB_D_FF_Float_58_70_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF58_70MultiplierStage1Output, mb_D_FF58_70MultiplierStage2Output);

    Multiplier_Float_58: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF58_70MultiplierStage2Output, flopocoMultiplier58WeightInput, Multiplier58_Output_70);

    MBRightSHR_Float_58_70: entity work.MBRightSHR(rtl)
    GENERIC MAP (43, NumberOfBits)
    PORT MAP (clk, rst, Multiplier58Weight, mbRightSHR58_70Output);

    MB_D_FF_Float_58_70_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR58_70Output, Multiplier58WeightOutput);

    InputIEEE_Float_58_70: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier58WeightOutput, flopocoMultiplier58WeightOutput);

    MB_D_FF_Float_58_70_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier58WeightOutput, flopocoMultiplier58WeightInput);

    MB_D_FF_Float_Multiplier18_61_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier8_Output_9, mb_D_FFMultiplier18_61_0Output);

    MB_D_FF_Float_61_73_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier18_61_0Output, mb_D_FF61_73MultiplierStage1Output);

    MB_D_FF_Float_61_73_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF61_73MultiplierStage1Output, mb_D_FF61_73MultiplierStage2Output);

    Multiplier_Float_61: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF61_73MultiplierStage2Output, flopocoMultiplier61WeightInput, Multiplier61_Output_73);

    MBRightSHR_Float_61_73: entity work.MBRightSHR(rtl)
    GENERIC MAP (43, NumberOfBits)
    PORT MAP (clk, rst, Multiplier61Weight, mbRightSHR61_73Output);

    MB_D_FF_Float_61_73_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR61_73Output, Multiplier61WeightOutput);

    InputIEEE_Float_61_73: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier61WeightOutput, flopocoMultiplier61WeightOutput);

    MB_D_FF_Float_61_73_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier61WeightOutput, flopocoMultiplier61WeightInput);

    MB_D_FF_Float_Adder17_Input1_12_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier61_Output_73, mb_D_FFAdder17_Input1_12_0Output);

    MB_D_FF_Float_12_74_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder17_Input1_12_0Output, mb_D_FF12_74AugendStage1Output);

    MB_D_FF_Float_12_74_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF12_74AugendStage1Output, mb_D_FF12_74AugendStage2Output);

    Adder_Float_12: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF12_74AugendStage2Output, mb_D_FF12_74AddendStage2Output, Adder12_Output_74);

    MB_D_FF_Float_Adder17_Input2_12_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier58_Output_70, mb_D_FFAdder17_Input2_12_0Output);

    MB_D_FF_Float_12_74_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder17_Input2_12_0Output, mb_D_FF12_74AddendStage1Output);

    MB_D_FF_Float_12_74_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF12_74AddendStage1Output, mb_D_FF12_74AddendStage2Output);

    MB_D_FF_Float_Multiplier16_Input1_62_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder12_Output_74, mb_D_FFMultiplier16_Input1_62_0Output);

    MB_D_FF_Float_62_75_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier16_Input1_62_0Output, mb_D_FF62_75MultiplicandStage1Output);

    MB_D_FF_Float_62_75_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF62_75MultiplicandStage1Output, mb_D_FF62_75MultiplicandStage2Output);

    Multiplier_Float_62: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF62_75MultiplicandStage2Output, mb_D_FF62_75MultiplierStage2Output, Multiplier62_Output_75);

    MB_D_FF_Float_Multiplier16_Input2_62_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier55_Output_67, mb_D_FFMultiplier16_Input2_62_0Output);

    MB_D_FF_Float_62_75_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier16_Input2_62_0Output, mb_D_FF62_75MultiplierStage1Output);

    MB_D_FF_Float_62_75_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF62_75MultiplierStage1Output, mb_D_FF62_75MultiplierStage2Output);

    MB_D_FF_Float_Multiplier15_63_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier62_Output_75, mb_D_FFMultiplier15_63_0Output);

    MB_D_FF_Float_63_76_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier15_63_0Output, mb_D_FF63_76MultiplierStage1Output);

    MB_D_FF_Float_63_76_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF63_76MultiplierStage1Output, mb_D_FF63_76MultiplierStage2Output);

    Multiplier_Float_63: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF63_76MultiplierStage2Output, flopocoMultiplier63WeightInput, Multiplier63_Output_76);

    MBRightSHR_Float_63_76: entity work.MBRightSHR(rtl)
    GENERIC MAP (82, NumberOfBits)
    PORT MAP (clk, rst, Multiplier63Weight, mbRightSHR63_76Output);

    MB_D_FF_Float_63_76_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR63_76Output, Multiplier63WeightOutput);

    InputIEEE_Float_63_76: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier63WeightOutput, flopocoMultiplier63WeightOutput);

    MB_D_FF_Float_63_76_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier63WeightOutput, flopocoMultiplier63WeightInput);

    MBRightSHR_Float_64_Input177: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits)
    PORT MAP (clk, rst, Multiplier64Weight, mbRightSHR64_Input1_77Output);

    MB_D_FF_Float_64_77_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR64_Input1_77Output, Multiplier64WeightOutput);

    InputIEEE_Float_64_77: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier64WeightOutput, flopocoMultiplier64WeightOutput);

    MB_D_FF_Float_64_77_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier64WeightOutput, flopocoMultiplier64WeightInput);

    Multiplier_Float_64: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier64WeightInput, mb_D_FF64_77MultiplierStage2Output, Multiplier64_Output_77);

    MBRightSHR_Float_64_Input2_77: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR64_Input2_77Input, mbRightSHR64_Input2_77Output);

    MB_D_FF_Float_64_77_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR64_Input2_77Output, mb_D_FF64_77MultiplierStage1Output);

    MB_D_FF_Float_64_77_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF64_77MultiplierStage1Output, mb_D_FF64_77MultiplierStage2Output);

    MBRightSHR_Float_65_Input178: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits)
    PORT MAP (clk, rst, Multiplier65Weight, mbRightSHR65_Input1_78Output);

    MB_D_FF_Float_65_78_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR65_Input1_78Output, Multiplier65WeightOutput);

    InputIEEE_Float_65_78: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier65WeightOutput, flopocoMultiplier65WeightOutput);

    MB_D_FF_Float_65_78_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier65WeightOutput, flopocoMultiplier65WeightInput);

    Multiplier_Float_65: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier65WeightInput, mb_D_FF65_78MultiplierStage2Output, Multiplier65_Output_78);

    MBRightSHR_Float_65_Input2_78: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR65_Input2_78Input, mbRightSHR65_Input2_78Output);

    MB_D_FF_Float_65_78_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR65_Input2_78Output, mb_D_FF65_78MultiplierStage1Output);

    MB_D_FF_Float_65_78_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF65_78MultiplierStage1Output, mb_D_FF65_78MultiplierStage2Output);

    MB_D_FF_Float_Adder18_Input1_13_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier65_Output_78, mb_D_FFAdder18_Input1_13_0Output);

    MB_D_FF_Float_13_79_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder18_Input1_13_0Output, mb_D_FF13_79AugendStage1Output);

    MB_D_FF_Float_13_79_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF13_79AugendStage1Output, mb_D_FF13_79AugendStage2Output);

    Adder_Float_13: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF13_79AugendStage2Output, mb_D_FF13_79AddendStage2Output, Adder13_Output_79);

    MB_D_FF_Float_Adder18_Input2_13_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier64_Output_77, mb_D_FFAdder18_Input2_13_0Output);

    MB_D_FF_Float_13_79_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder18_Input2_13_0Output, mb_D_FF13_79AddendStage1Output);

    MB_D_FF_Float_13_79_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF13_79AddendStage1Output, mb_D_FF13_79AddendStage2Output);

    MB_D_FF_Float_Multiplier17_66_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder13_Output_79, mb_D_FFMultiplier17_66_0Output);

    MB_D_FF_Float_66_80_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier17_66_0Output, mb_D_FF66_80MultiplierStage1Output);

    MB_D_FF_Float_66_80_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF66_80MultiplierStage1Output, mb_D_FF66_80MultiplierStage2Output);

    Multiplier_Float_66: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF66_80MultiplierStage2Output, mb_D_FF66_80MultiplicandStage2Output, Multiplier66_Output_80);

    MBRightSHR_Float_66_80: entity work.MBRightSHR(rtl)
    GENERIC MAP (50, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR66_80Input, mbRightSHR66_80Output);

    MB_D_FF_Float_66_80_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR66_80Output, mb_D_FF66_80MultiplicandStage1Output);

    MB_D_FF_Float_66_80_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF66_80MultiplicandStage1Output, mb_D_FF66_80MultiplicandStage2Output);

    MB_D_FF_Float_Multiplier18_69_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier16_Output_19, mb_D_FFMultiplier18_69_0Output);

    MB_D_FF_Float_69_83_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier18_69_0Output, mb_D_FF69_83MultiplierStage1Output);

    MB_D_FF_Float_69_83_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF69_83MultiplierStage1Output, mb_D_FF69_83MultiplierStage2Output);

    Multiplier_Float_69: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF69_83MultiplierStage2Output, flopocoMultiplier69WeightInput, Multiplier69_Output_83);

    MBRightSHR_Float_69_83: entity work.MBRightSHR(rtl)
    GENERIC MAP (43, NumberOfBits)
    PORT MAP (clk, rst, Multiplier69Weight, mbRightSHR69_83Output);

    MB_D_FF_Float_69_83_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR69_83Output, Multiplier69WeightOutput);

    InputIEEE_Float_69_83: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier69WeightOutput, flopocoMultiplier69WeightOutput);

    MB_D_FF_Float_69_83_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier69WeightOutput, flopocoMultiplier69WeightInput);

    MB_D_FF_Float_Multiplier18_72_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier19_Output_22, mb_D_FFMultiplier18_72_0Output);

    MB_D_FF_Float_72_86_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier18_72_0Output, mb_D_FF72_86MultiplierStage1Output);

    MB_D_FF_Float_72_86_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF72_86MultiplierStage1Output, mb_D_FF72_86MultiplierStage2Output);

    Multiplier_Float_72: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF72_86MultiplierStage2Output, flopocoMultiplier72WeightInput, Multiplier72_Output_86);

    MBRightSHR_Float_72_86: entity work.MBRightSHR(rtl)
    GENERIC MAP (43, NumberOfBits)
    PORT MAP (clk, rst, Multiplier72Weight, mbRightSHR72_86Output);

    MB_D_FF_Float_72_86_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR72_86Output, Multiplier72WeightOutput);

    InputIEEE_Float_72_86: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier72WeightOutput, flopocoMultiplier72WeightOutput);

    MB_D_FF_Float_72_86_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier72WeightOutput, flopocoMultiplier72WeightInput);

    MB_D_FF_Float_Adder17_Input1_14_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier72_Output_86, mb_D_FFAdder17_Input1_14_0Output);

    MB_D_FF_Float_14_87_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder17_Input1_14_0Output, mb_D_FF14_87AugendStage1Output);

    MB_D_FF_Float_14_87_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF14_87AugendStage1Output, mb_D_FF14_87AugendStage2Output);

    Adder_Float_14: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF14_87AugendStage2Output, mb_D_FF14_87AddendStage2Output, Adder14_Output_87);

    MB_D_FF_Float_Adder17_Input2_14_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier69_Output_83, mb_D_FFAdder17_Input2_14_0Output);

    MB_D_FF_Float_14_87_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder17_Input2_14_0Output, mb_D_FF14_87AddendStage1Output);

    MB_D_FF_Float_14_87_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF14_87AddendStage1Output, mb_D_FF14_87AddendStage2Output);

    MB_D_FF_Float_Multiplier16_Input1_73_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder14_Output_87, mb_D_FFMultiplier16_Input1_73_0Output);

    MB_D_FF_Float_73_88_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier16_Input1_73_0Output, mb_D_FF73_88MultiplicandStage1Output);

    MB_D_FF_Float_73_88_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF73_88MultiplicandStage1Output, mb_D_FF73_88MultiplicandStage2Output);

    Multiplier_Float_73: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF73_88MultiplicandStage2Output, mb_D_FF73_88MultiplierStage2Output, Multiplier73_Output_88);

    MB_D_FF_Float_Multiplier16_Input2_73_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier66_Output_80, mb_D_FFMultiplier16_Input2_73_0Output);

    MB_D_FF_Float_73_88_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier16_Input2_73_0Output, mb_D_FF73_88MultiplierStage1Output);

    MB_D_FF_Float_73_88_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF73_88MultiplierStage1Output, mb_D_FF73_88MultiplierStage2Output);

    MB_D_FF_Float_Multiplier15_74_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier73_Output_88, mb_D_FFMultiplier15_74_0Output);

    MB_D_FF_Float_74_89_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier15_74_0Output, mb_D_FF74_89MultiplierStage1Output);

    MB_D_FF_Float_74_89_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF74_89MultiplierStage1Output, mb_D_FF74_89MultiplierStage2Output);

    Multiplier_Float_74: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF74_89MultiplierStage2Output, flopocoMultiplier74WeightInput, Multiplier74_Output_89);

    MBRightSHR_Float_74_89: entity work.MBRightSHR(rtl)
    GENERIC MAP (82, NumberOfBits)
    PORT MAP (clk, rst, Multiplier74Weight, mbRightSHR74_89Output);

    MB_D_FF_Float_74_89_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR74_89Output, Multiplier74WeightOutput);

    InputIEEE_Float_74_89: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier74WeightOutput, flopocoMultiplier74WeightOutput);

    MB_D_FF_Float_74_89_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier74WeightOutput, flopocoMultiplier74WeightInput);

    MB_D_FF_Float_Adder14_Input1_15_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier74_Output_89, mb_D_FFAdder14_Input1_15_0Output);

    MB_D_FF_Float_15_90_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder14_Input1_15_0Output, mb_D_FF15_90AugendStage1Output);

    MB_D_FF_Float_15_90_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF15_90AugendStage1Output, mb_D_FF15_90AugendStage2Output);

    Adder_Float_15: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF15_90AugendStage2Output, mb_D_FF15_90AddendStage2Output, Adder15_Output_90);

    MB_D_FF_Float_Adder14_Input2_15_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier63_Output_76, mb_D_FFAdder14_Input2_15_0Output);

    MB_D_FF_Float_15_90_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder14_Input2_15_0Output, mb_D_FF15_90AddendStage1Output);

    MB_D_FF_Float_15_90_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF15_90AddendStage1Output, mb_D_FF15_90AddendStage2Output);

    MB_D_FF_Float_Multiplier13_Input1_75_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder15_Output_90, mb_D_FFMultiplier13_Input1_75_0Output);

    MB_D_FF_Float_75_91_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier13_Input1_75_0Output, mb_D_FF75_91MultiplicandStage1Output);

    MB_D_FF_Float_75_91_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF75_91MultiplicandStage1Output, mb_D_FF75_91MultiplicandStage2Output);

    Multiplier_Float_75: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF75_91MultiplicandStage2Output, mb_D_FF75_91MultiplierStage2Output, Multiplier75_Output_91);

    MB_D_FF_Float_Multiplier13_Input2_75_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier0_Output_0, mb_D_FFMultiplier13_Input2_75_0Output);

    MB_D_FF_Float_75_91_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier13_Input2_75_0Output, mb_D_FF75_91MultiplierStage1Output);

    MB_D_FF_Float_75_91_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF75_91MultiplierStage1Output, mb_D_FF75_91MultiplierStage2Output);

    MB_D_FF_Float_Multiplier12_76_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier75_Output_91, mb_D_FFMultiplier12_76_0Output);

    MB_D_FF_Float_76_92_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier12_76_0Output, mb_D_FF76_92MultiplierStage1Output);

    MB_D_FF_Float_76_92_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF76_92MultiplierStage1Output, mb_D_FF76_92MultiplierStage2Output);

    Multiplier_Float_76: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF76_92MultiplierStage2Output, flopocoMultiplier76WeightInput, Multiplier76_Output_92);

    MBRightSHR_Float_76_92: entity work.MBRightSHR(rtl)
    GENERIC MAP (121, NumberOfBits)
    PORT MAP (clk, rst, Multiplier76Weight, mbRightSHR76_92Output);

    MB_D_FF_Float_76_92_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR76_92Output, Multiplier76WeightOutput);

    InputIEEE_Float_76_92: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier76WeightOutput, flopocoMultiplier76WeightOutput);

    MB_D_FF_Float_76_92_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier76WeightOutput, flopocoMultiplier76WeightInput);

    MBRightSHR_Float_78_Input194: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits)
    PORT MAP (clk, rst, Multiplier78Weight, mbRightSHR78_Input1_94Output);

    MB_D_FF_Float_78_94_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR78_Input1_94Output, Multiplier78WeightOutput);

    InputIEEE_Float_78_94: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier78WeightOutput, flopocoMultiplier78WeightOutput);

    MB_D_FF_Float_78_94_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier78WeightOutput, flopocoMultiplier78WeightInput);

    Multiplier_Float_78: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier78WeightInput, mb_D_FF78_94MultiplierStage2Output, Multiplier78_Output_94);

    MBRightSHR_Float_78_Input2_94: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR78_Input2_94Input, mbRightSHR78_Input2_94Output);

    MB_D_FF_Float_78_94_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR78_Input2_94Output, mb_D_FF78_94MultiplierStage1Output);

    MB_D_FF_Float_78_94_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF78_94MultiplierStage1Output, mb_D_FF78_94MultiplierStage2Output);

    MBRightSHR_Float_79_Input195: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits)
    PORT MAP (clk, rst, Multiplier79Weight, mbRightSHR79_Input1_95Output);

    MB_D_FF_Float_79_95_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR79_Input1_95Output, Multiplier79WeightOutput);

    InputIEEE_Float_79_95: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier79WeightOutput, flopocoMultiplier79WeightOutput);

    MB_D_FF_Float_79_95_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier79WeightOutput, flopocoMultiplier79WeightInput);

    Multiplier_Float_79: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier79WeightInput, mb_D_FF79_95MultiplierStage2Output, Multiplier79_Output_95);

    MBRightSHR_Float_79_Input2_95: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR79_Input2_95Input, mbRightSHR79_Input2_95Output);

    MB_D_FF_Float_79_95_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR79_Input2_95Output, mb_D_FF79_95MultiplierStage1Output);

    MB_D_FF_Float_79_95_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF79_95MultiplierStage1Output, mb_D_FF79_95MultiplierStage2Output);

    MB_D_FF_Float_Adder18_Input1_16_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier79_Output_95, mb_D_FFAdder18_Input1_16_0Output);

    MB_D_FF_Float_16_96_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder18_Input1_16_0Output, mb_D_FF16_96AugendStage1Output);

    MB_D_FF_Float_16_96_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF16_96AugendStage1Output, mb_D_FF16_96AugendStage2Output);

    Adder_Float_16: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF16_96AugendStage2Output, mb_D_FF16_96AddendStage2Output, Adder16_Output_96);

    MB_D_FF_Float_Adder18_Input2_16_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier78_Output_94, mb_D_FFAdder18_Input2_16_0Output);

    MB_D_FF_Float_16_96_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder18_Input2_16_0Output, mb_D_FF16_96AddendStage1Output);

    MB_D_FF_Float_16_96_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF16_96AddendStage1Output, mb_D_FF16_96AddendStage2Output);

    MB_D_FF_Float_Multiplier17_80_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder16_Output_96, mb_D_FFMultiplier17_80_0Output);

    MB_D_FF_Float_80_97_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier17_80_0Output, mb_D_FF80_97MultiplierStage1Output);

    MB_D_FF_Float_80_97_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF80_97MultiplierStage1Output, mb_D_FF80_97MultiplierStage2Output);

    Multiplier_Float_80: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF80_97MultiplierStage2Output, mb_D_FF80_97MultiplicandStage2Output, Multiplier80_Output_97);

    MBRightSHR_Float_80_97: entity work.MBRightSHR(rtl)
    GENERIC MAP (50, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR80_97Input, mbRightSHR80_97Output);

    MB_D_FF_Float_80_97_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR80_97Output, mb_D_FF80_97MultiplicandStage1Output);

    MB_D_FF_Float_80_97_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF80_97MultiplicandStage1Output, mb_D_FF80_97MultiplicandStage2Output);

    MB_D_FF_Float_Multiplier18_83_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier30_Output_36, mb_D_FFMultiplier18_83_0Output);

    MB_D_FF_Float_83_100_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier18_83_0Output, mb_D_FF83_100MultiplierStage1Output);

    MB_D_FF_Float_83_100_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF83_100MultiplierStage1Output, mb_D_FF83_100MultiplierStage2Output);

    Multiplier_Float_83: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF83_100MultiplierStage2Output, flopocoMultiplier83WeightInput, Multiplier83_Output_100);

    MBRightSHR_Float_83_100: entity work.MBRightSHR(rtl)
    GENERIC MAP (43, NumberOfBits)
    PORT MAP (clk, rst, Multiplier83Weight, mbRightSHR83_100Output);

    MB_D_FF_Float_83_100_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR83_100Output, Multiplier83WeightOutput);

    InputIEEE_Float_83_100: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier83WeightOutput, flopocoMultiplier83WeightOutput);

    MB_D_FF_Float_83_100_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier83WeightOutput, flopocoMultiplier83WeightInput);

    MB_D_FF_Float_Multiplier18_86_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier33_Output_39, mb_D_FFMultiplier18_86_0Output);

    MB_D_FF_Float_86_103_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier18_86_0Output, mb_D_FF86_103MultiplierStage1Output);

    MB_D_FF_Float_86_103_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF86_103MultiplierStage1Output, mb_D_FF86_103MultiplierStage2Output);

    Multiplier_Float_86: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF86_103MultiplierStage2Output, flopocoMultiplier86WeightInput, Multiplier86_Output_103);

    MBRightSHR_Float_86_103: entity work.MBRightSHR(rtl)
    GENERIC MAP (43, NumberOfBits)
    PORT MAP (clk, rst, Multiplier86Weight, mbRightSHR86_103Output);

    MB_D_FF_Float_86_103_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR86_103Output, Multiplier86WeightOutput);

    InputIEEE_Float_86_103: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier86WeightOutput, flopocoMultiplier86WeightOutput);

    MB_D_FF_Float_86_103_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier86WeightOutput, flopocoMultiplier86WeightInput);

    MB_D_FF_Float_Adder17_Input1_17_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier86_Output_103, mb_D_FFAdder17_Input1_17_0Output);

    MB_D_FF_Float_17_104_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder17_Input1_17_0Output, mb_D_FF17_104AugendStage1Output);

    MB_D_FF_Float_17_104_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF17_104AugendStage1Output, mb_D_FF17_104AugendStage2Output);

    Adder_Float_17: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF17_104AugendStage2Output, mb_D_FF17_104AddendStage2Output, Adder17_Output_104);

    MB_D_FF_Float_Adder17_Input2_17_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier83_Output_100, mb_D_FFAdder17_Input2_17_0Output);

    MB_D_FF_Float_17_104_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder17_Input2_17_0Output, mb_D_FF17_104AddendStage1Output);

    MB_D_FF_Float_17_104_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF17_104AddendStage1Output, mb_D_FF17_104AddendStage2Output);

    MB_D_FF_Float_Multiplier16_Input1_87_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder17_Output_104, mb_D_FFMultiplier16_Input1_87_0Output);

    MB_D_FF_Float_87_105_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier16_Input1_87_0Output, mb_D_FF87_105MultiplicandStage1Output);

    MB_D_FF_Float_87_105_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF87_105MultiplicandStage1Output, mb_D_FF87_105MultiplicandStage2Output);

    Multiplier_Float_87: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF87_105MultiplicandStage2Output, mb_D_FF87_105MultiplierStage2Output, Multiplier87_Output_105);

    MB_D_FF_Float_Multiplier16_Input2_87_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier80_Output_97, mb_D_FFMultiplier16_Input2_87_0Output);

    MB_D_FF_Float_87_105_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier16_Input2_87_0Output, mb_D_FF87_105MultiplierStage1Output);

    MB_D_FF_Float_87_105_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF87_105MultiplierStage1Output, mb_D_FF87_105MultiplierStage2Output);

    MB_D_FF_Float_Multiplier15_88_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier87_Output_105, mb_D_FFMultiplier15_88_0Output);

    MB_D_FF_Float_88_106_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier15_88_0Output, mb_D_FF88_106MultiplierStage1Output);

    MB_D_FF_Float_88_106_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF88_106MultiplierStage1Output, mb_D_FF88_106MultiplierStage2Output);

    Multiplier_Float_88: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF88_106MultiplierStage2Output, flopocoMultiplier88WeightInput, Multiplier88_Output_106);

    MBRightSHR_Float_88_106: entity work.MBRightSHR(rtl)
    GENERIC MAP (82, NumberOfBits)
    PORT MAP (clk, rst, Multiplier88Weight, mbRightSHR88_106Output);

    MB_D_FF_Float_88_106_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR88_106Output, Multiplier88WeightOutput);

    InputIEEE_Float_88_106: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier88WeightOutput, flopocoMultiplier88WeightOutput);

    MB_D_FF_Float_88_106_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier88WeightOutput, flopocoMultiplier88WeightInput);

    MBRightSHR_Float_89_Input1107: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits)
    PORT MAP (clk, rst, Multiplier89Weight, mbRightSHR89_Input1_107Output);

    MB_D_FF_Float_89_107_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR89_Input1_107Output, Multiplier89WeightOutput);

    InputIEEE_Float_89_107: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier89WeightOutput, flopocoMultiplier89WeightOutput);

    MB_D_FF_Float_89_107_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier89WeightOutput, flopocoMultiplier89WeightInput);

    Multiplier_Float_89: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier89WeightInput, mb_D_FF89_107MultiplierStage2Output, Multiplier89_Output_107);

    MBRightSHR_Float_89_Input2_107: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR89_Input2_107Input, mbRightSHR89_Input2_107Output);

    MB_D_FF_Float_89_107_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR89_Input2_107Output, mb_D_FF89_107MultiplierStage1Output);

    MB_D_FF_Float_89_107_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF89_107MultiplierStage1Output, mb_D_FF89_107MultiplierStage2Output);

    MBRightSHR_Float_90_Input1108: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits)
    PORT MAP (clk, rst, Multiplier90Weight, mbRightSHR90_Input1_108Output);

    MB_D_FF_Float_90_108_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR90_Input1_108Output, Multiplier90WeightOutput);

    InputIEEE_Float_90_108: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier90WeightOutput, flopocoMultiplier90WeightOutput);

    MB_D_FF_Float_90_108_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier90WeightOutput, flopocoMultiplier90WeightInput);

    Multiplier_Float_90: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier90WeightInput, mb_D_FF90_108MultiplierStage2Output, Multiplier90_Output_108);

    MBRightSHR_Float_90_Input2_108: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR90_Input2_108Input, mbRightSHR90_Input2_108Output);

    MB_D_FF_Float_90_108_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR90_Input2_108Output, mb_D_FF90_108MultiplierStage1Output);

    MB_D_FF_Float_90_108_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF90_108MultiplierStage1Output, mb_D_FF90_108MultiplierStage2Output);

    MB_D_FF_Float_Adder18_Input1_18_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier90_Output_108, mb_D_FFAdder18_Input1_18_0Output);

    MB_D_FF_Float_18_109_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder18_Input1_18_0Output, mb_D_FF18_109AugendStage1Output);

    MB_D_FF_Float_18_109_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF18_109AugendStage1Output, mb_D_FF18_109AugendStage2Output);

    Adder_Float_18: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF18_109AugendStage2Output, mb_D_FF18_109AddendStage2Output, Adder18_Output_109);

    MB_D_FF_Float_Adder18_Input2_18_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier89_Output_107, mb_D_FFAdder18_Input2_18_0Output);

    MB_D_FF_Float_18_109_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder18_Input2_18_0Output, mb_D_FF18_109AddendStage1Output);

    MB_D_FF_Float_18_109_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF18_109AddendStage1Output, mb_D_FF18_109AddendStage2Output);

    MB_D_FF_Float_Multiplier17_91_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder18_Output_109, mb_D_FFMultiplier17_91_0Output);

    MB_D_FF_Float_91_110_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier17_91_0Output, mb_D_FF91_110MultiplierStage1Output);

    MB_D_FF_Float_91_110_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF91_110MultiplierStage1Output, mb_D_FF91_110MultiplierStage2Output);

    Multiplier_Float_91: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF91_110MultiplierStage2Output, mb_D_FF91_110MultiplicandStage2Output, Multiplier91_Output_110);

    MBRightSHR_Float_91_110: entity work.MBRightSHR(rtl)
    GENERIC MAP (50, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR91_110Input, mbRightSHR91_110Output);

    MB_D_FF_Float_91_110_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR91_110Output, mb_D_FF91_110MultiplicandStage1Output);

    MB_D_FF_Float_91_110_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF91_110MultiplicandStage1Output, mb_D_FF91_110MultiplicandStage2Output);

    MB_D_FF_Float_Multiplier18_94_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier41_Output_49, mb_D_FFMultiplier18_94_0Output);

    MB_D_FF_Float_94_113_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier18_94_0Output, mb_D_FF94_113MultiplierStage1Output);

    MB_D_FF_Float_94_113_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF94_113MultiplierStage1Output, mb_D_FF94_113MultiplierStage2Output);

    Multiplier_Float_94: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF94_113MultiplierStage2Output, flopocoMultiplier94WeightInput, Multiplier94_Output_113);

    MBRightSHR_Float_94_113: entity work.MBRightSHR(rtl)
    GENERIC MAP (43, NumberOfBits)
    PORT MAP (clk, rst, Multiplier94Weight, mbRightSHR94_113Output);

    MB_D_FF_Float_94_113_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR94_113Output, Multiplier94WeightOutput);

    InputIEEE_Float_94_113: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier94WeightOutput, flopocoMultiplier94WeightOutput);

    MB_D_FF_Float_94_113_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier94WeightOutput, flopocoMultiplier94WeightInput);

    MB_D_FF_Float_Multiplier18_97_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier44_Output_52, mb_D_FFMultiplier18_97_0Output);

    MB_D_FF_Float_97_116_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier18_97_0Output, mb_D_FF97_116MultiplierStage1Output);

    MB_D_FF_Float_97_116_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF97_116MultiplierStage1Output, mb_D_FF97_116MultiplierStage2Output);

    Multiplier_Float_97: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF97_116MultiplierStage2Output, flopocoMultiplier97WeightInput, Multiplier97_Output_116);

    MBRightSHR_Float_97_116: entity work.MBRightSHR(rtl)
    GENERIC MAP (43, NumberOfBits)
    PORT MAP (clk, rst, Multiplier97Weight, mbRightSHR97_116Output);

    MB_D_FF_Float_97_116_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR97_116Output, Multiplier97WeightOutput);

    InputIEEE_Float_97_116: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier97WeightOutput, flopocoMultiplier97WeightOutput);

    MB_D_FF_Float_97_116_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier97WeightOutput, flopocoMultiplier97WeightInput);

    MB_D_FF_Float_Adder17_Input1_19_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier97_Output_116, mb_D_FFAdder17_Input1_19_0Output);

    MB_D_FF_Float_19_117_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder17_Input1_19_0Output, mb_D_FF19_117AugendStage1Output);

    MB_D_FF_Float_19_117_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF19_117AugendStage1Output, mb_D_FF19_117AugendStage2Output);

    Adder_Float_19: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF19_117AugendStage2Output, mb_D_FF19_117AddendStage2Output, Adder19_Output_117);

    MB_D_FF_Float_Adder17_Input2_19_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier94_Output_113, mb_D_FFAdder17_Input2_19_0Output);

    MB_D_FF_Float_19_117_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder17_Input2_19_0Output, mb_D_FF19_117AddendStage1Output);

    MB_D_FF_Float_19_117_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF19_117AddendStage1Output, mb_D_FF19_117AddendStage2Output);

    MB_D_FF_Float_Multiplier16_Input1_98_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder19_Output_117, mb_D_FFMultiplier16_Input1_98_0Output);

    MB_D_FF_Float_98_118_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier16_Input1_98_0Output, mb_D_FF98_118MultiplicandStage1Output);

    MB_D_FF_Float_98_118_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF98_118MultiplicandStage1Output, mb_D_FF98_118MultiplicandStage2Output);

    Multiplier_Float_98: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF98_118MultiplicandStage2Output, mb_D_FF98_118MultiplierStage2Output, Multiplier98_Output_118);

    MB_D_FF_Float_Multiplier16_Input2_98_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier91_Output_110, mb_D_FFMultiplier16_Input2_98_0Output);

    MB_D_FF_Float_98_118_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier16_Input2_98_0Output, mb_D_FF98_118MultiplierStage1Output);

    MB_D_FF_Float_98_118_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF98_118MultiplierStage1Output, mb_D_FF98_118MultiplierStage2Output);

    MB_D_FF_Float_Multiplier15_99_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier98_Output_118, mb_D_FFMultiplier15_99_0Output);

    MB_D_FF_Float_99_119_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier15_99_0Output, mb_D_FF99_119MultiplierStage1Output);

    MB_D_FF_Float_99_119_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF99_119MultiplierStage1Output, mb_D_FF99_119MultiplierStage2Output);

    Multiplier_Float_99: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF99_119MultiplierStage2Output, flopocoMultiplier99WeightInput, Multiplier99_Output_119);

    MBRightSHR_Float_99_119: entity work.MBRightSHR(rtl)
    GENERIC MAP (82, NumberOfBits)
    PORT MAP (clk, rst, Multiplier99Weight, mbRightSHR99_119Output);

    MB_D_FF_Float_99_119_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR99_119Output, Multiplier99WeightOutput);

    InputIEEE_Float_99_119: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier99WeightOutput, flopocoMultiplier99WeightOutput);

    MB_D_FF_Float_99_119_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier99WeightOutput, flopocoMultiplier99WeightInput);

    MB_D_FF_Float_Adder14_Input1_20_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier99_Output_119, mb_D_FFAdder14_Input1_20_0Output);

    MB_D_FF_Float_20_120_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder14_Input1_20_0Output, mb_D_FF20_120AugendStage1Output);

    MB_D_FF_Float_20_120_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF20_120AugendStage1Output, mb_D_FF20_120AugendStage2Output);

    Adder_Float_20: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF20_120AugendStage2Output, mb_D_FF20_120AddendStage2Output, Adder20_Output_120);

    MB_D_FF_Float_Adder14_Input2_20_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier88_Output_106, mb_D_FFAdder14_Input2_20_0Output);

    MB_D_FF_Float_20_120_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder14_Input2_20_0Output, mb_D_FF20_120AddendStage1Output);

    MB_D_FF_Float_20_120_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF20_120AddendStage1Output, mb_D_FF20_120AddendStage2Output);

    MB_D_FF_Float_Multiplier13_Input1_100_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder20_Output_120, mb_D_FFMultiplier13_Input1_100_0Output);

    MB_D_FF_Float_100_121_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier13_Input1_100_0Output, mb_D_FF100_121MultiplicandStage1Output);

    MB_D_FF_Float_100_121_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF100_121MultiplicandStage1Output, mb_D_FF100_121MultiplicandStage2Output);

    Multiplier_Float_100: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF100_121MultiplicandStage2Output, mb_D_FF100_121MultiplierStage2Output, Multiplier100_Output_121);

    MB_D_FF_Float_Multiplier13_Input2_100_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier25_Output_30, mb_D_FFMultiplier13_Input2_100_0Output);

    MB_D_FF_Float_100_121_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier13_Input2_100_0Output, mb_D_FF100_121MultiplierStage1Output);

    MB_D_FF_Float_100_121_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF100_121MultiplierStage1Output, mb_D_FF100_121MultiplierStage2Output);

    MB_D_FF_Float_Multiplier12_101_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier100_Output_121, mb_D_FFMultiplier12_101_0Output);

    MB_D_FF_Float_101_122_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier12_101_0Output, mb_D_FF101_122MultiplierStage1Output);

    MB_D_FF_Float_101_122_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF101_122MultiplierStage1Output, mb_D_FF101_122MultiplierStage2Output);

    Multiplier_Float_101: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF101_122MultiplierStage2Output, flopocoMultiplier101WeightInput, Multiplier101_Output_122);

    MBRightSHR_Float_101_122: entity work.MBRightSHR(rtl)
    GENERIC MAP (121, NumberOfBits)
    PORT MAP (clk, rst, Multiplier101Weight, mbRightSHR101_122Output);

    MB_D_FF_Float_101_122_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR101_122Output, Multiplier101WeightOutput);

    InputIEEE_Float_101_122: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier101WeightOutput, flopocoMultiplier101WeightOutput);

    MB_D_FF_Float_101_122_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier101WeightOutput, flopocoMultiplier101WeightInput);

    MB_D_FF_Float_Adder11_Input1_21_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier101_Output_122, mb_D_FFAdder11_Input1_21_0Output);

    MB_D_FF_Float_21_123_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder11_Input1_21_0Output, mb_D_FF21_123AugendStage1Output);

    MB_D_FF_Float_21_123_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF21_123AugendStage1Output, mb_D_FF21_123AugendStage2Output);

    Adder_Float_21: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF21_123AugendStage2Output, mb_D_FF21_123AddendStage2Output, Adder21_Output_123);

    MB_D_FF_Float_Adder11_Input2_21_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier76_Output_92, mb_D_FFAdder11_Input2_21_0Output);

    MB_D_FF_Float_21_123_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder11_Input2_21_0Output, mb_D_FF21_123AddendStage1Output);

    MB_D_FF_Float_21_123_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF21_123AddendStage1Output, mb_D_FF21_123AddendStage2Output);

    MB_D_FF_Float_Multiplier10_102_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder21_Output_123, mb_D_FFMultiplier10_102_0Output);

    MB_D_FF_Float_102_124_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier10_102_0Output, mb_D_FF102_124MultiplierStage1Output);

    MB_D_FF_Float_102_124_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF102_124MultiplierStage1Output, mb_D_FF102_124MultiplierStage2Output);

    Multiplier_Float_102: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF102_124MultiplierStage2Output, mb_D_FF102_124MultiplicandStage2Output, Multiplier102_Output_124);

    MBRightSHR_Float_102_124: entity work.MBRightSHR(rtl)
    GENERIC MAP (135, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR102_124Input, mbRightSHR102_124Output);

    MB_D_FF_Float_102_124_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR102_124Output, mb_D_FF102_124MultiplicandStage1Output);

    MB_D_FF_Float_102_124_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF102_124MultiplicandStage1Output, mb_D_FF102_124MultiplicandStage2Output);

    MB_D_FF_Float_Multiplier9_103_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier102_Output_124, mb_D_FFMultiplier9_103_0Output);

    MB_D_FF_Float_103_125_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier9_103_0Output, mb_D_FF103_125MultiplierStage1Output);

    MB_D_FF_Float_103_125_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF103_125MultiplierStage1Output, mb_D_FF103_125MultiplierStage2Output);

    Multiplier_Float_103: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF103_125MultiplierStage2Output, flopocoMultiplier103WeightInput, Multiplier103_Output_125);

    MBRightSHR_Float_103_125: entity work.MBRightSHR(rtl)
    GENERIC MAP (160, NumberOfBits)
    PORT MAP (clk, rst, Multiplier103Weight, mbRightSHR103_125Output);

    MB_D_FF_Float_103_125_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR103_125Output, Multiplier103WeightOutput);

    InputIEEE_Float_103_125: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier103WeightOutput, flopocoMultiplier103WeightOutput);

    MB_D_FF_Float_103_125_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier103WeightOutput, flopocoMultiplier103WeightInput);

    MB_D_FF_Float_Adder8_Input1_22_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier103_Output_125, mb_D_FFAdder8_Input1_22_0Output);

    MB_D_FF_Float_22_126_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder8_Input1_22_0Output, mb_D_FF22_126AugendStage1Output);

    MB_D_FF_Float_22_126_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF22_126AugendStage1Output, mb_D_FF22_126AugendStage2Output);

    Adder_Float_22: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF22_126AugendStage2Output, mb_D_FF22_126AddendStage2Output, Adder22_Output_126);

    MB_D_FF_Float_Adder8_Input2_22_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier51_Output_62, mb_D_FFAdder8_Input2_22_0Output);

    MB_D_FF_Float_22_126_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder8_Input2_22_0Output, mb_D_FF22_126AddendStage1Output);

    MB_D_FF_Float_22_126_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF22_126AddendStage1Output, mb_D_FF22_126AddendStage2Output);

    MB_D_FF_Float_Multiplier7_104_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder22_Output_126, mb_D_FFMultiplier7_104_0Output);

    MB_D_FF_Float_104_127_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier7_104_0Output, mb_D_FF104_127MultiplierStage1Output);

    MB_D_FF_Float_104_127_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF104_127MultiplierStage1Output, mb_D_FF104_127MultiplierStage2Output);

    Multiplier_Float_104: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF104_127MultiplierStage2Output, mb_D_FF104_127MultiplicandStage2Output, Multiplier104_Output_127);

    MBRightSHR_Float_104_127: entity work.MBRightSHR(rtl)
    GENERIC MAP (174, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR104_127Input, mbRightSHR104_127Output);

    MB_D_FF_Float_104_127_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR104_127Output, mb_D_FF104_127MultiplicandStage1Output);

    MB_D_FF_Float_104_127_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF104_127MultiplicandStage1Output, mb_D_FF104_127MultiplicandStage2Output);

    MBRightSHR_Float_105_128: entity work.MBRightSHR(rtl)
    GENERIC MAP (4, NumberOfBits)
    PORT MAP (clk, rst, Multiplier105Weight, mbRightSHR105_128Output);

    MB_D_FF_Float_105_128_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR105_128Output, Multiplier105WeightOutput);

    InputIEEE_Float_105_128: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier105WeightOutput, flopocoMultiplier105WeightOutput);

    MB_D_FF_Float_105_128_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier105WeightOutput, flopocoMultiplier105WeightInput);

    Multiplier_Float_105: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier105WeightInput, mb_D_FF105_128MultiplierStage2Output, Multiplier105_Output_128);

    MB_D_FF_Float_Multiplier21_105_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier21_105_0Input, mb_D_FFMultiplier21_105_0Output);

    MB_D_FF_Float_105_128_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier21_105_0Output, mb_D_FF105_128MultiplierStage1Output);

    MB_D_FF_Float_105_128_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF105_128MultiplierStage1Output, mb_D_FF105_128MultiplierStage2Output);

    MBRightSHR_Float_106_129: entity work.MBRightSHR(rtl)
    GENERIC MAP (4, NumberOfBits)
    PORT MAP (clk, rst, Multiplier106Weight, mbRightSHR106_129Output);

    MB_D_FF_Float_106_129_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR106_129Output, Multiplier106WeightOutput);

    InputIEEE_Float_106_129: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier106WeightOutput, flopocoMultiplier106WeightOutput);

    MB_D_FF_Float_106_129_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier106WeightOutput, flopocoMultiplier106WeightInput);

    Multiplier_Float_106: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier106WeightInput, mb_D_FF106_129MultiplierStage2Output, Multiplier106_Output_129);

    MB_D_FF_Float_Multiplier21_106_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier21_106_0Input, mb_D_FFMultiplier21_106_0Output);

    MB_D_FF_Float_106_129_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier21_106_0Output, mb_D_FF106_129MultiplierStage1Output);

    MB_D_FF_Float_106_129_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF106_129MultiplierStage1Output, mb_D_FF106_129MultiplierStage2Output);

    MB_D_FF_Float_Adder20_Input1_23_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier106_Output_129, mb_D_FFAdder20_Input1_23_0Output);

    MB_D_FF_Float_23_130_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder20_Input1_23_0Output, mb_D_FF23_130AugendStage1Output);

    MB_D_FF_Float_23_130_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF23_130AugendStage1Output, mb_D_FF23_130AugendStage2Output);

    Adder_Float_23: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF23_130AugendStage2Output, mb_D_FF23_130AddendStage2Output, Adder23_Output_130);

    MB_D_FF_Float_Adder20_Input2_23_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier105_Output_128, mb_D_FFAdder20_Input2_23_0Output);

    MB_D_FF_Float_23_130_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder20_Input2_23_0Output, mb_D_FF23_130AddendStage1Output);

    MB_D_FF_Float_23_130_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF23_130AddendStage1Output, mb_D_FF23_130AddendStage2Output);

    MB_D_FF_Float_Multiplier19_107_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder23_Output_130, mb_D_FFMultiplier19_107_0Output);

    MB_D_FF_Float_107_131_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier19_107_0Output, mb_D_FF107_131MultiplierStage1Output);

    MB_D_FF_Float_107_131_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF107_131MultiplierStage1Output, mb_D_FF107_131MultiplierStage2Output);

    Multiplier_Float_107: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF107_131MultiplierStage2Output, mb_D_FF107_131MultiplicandStage2Output, Multiplier107_Output_131);

    MBRightSHR_Float_107_131: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR107_131Input, mbRightSHR107_131Output);

    MB_D_FF_Float_107_131_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR107_131Output, mb_D_FF107_131MultiplicandStage1Output);

    MB_D_FF_Float_107_131_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF107_131MultiplicandStage1Output, mb_D_FF107_131MultiplicandStage2Output);

    MB_D_FF_Float_Multiplier18_108_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier107_Output_131, mb_D_FFMultiplier18_108_0Output);

    MB_D_FF_Float_108_132_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier18_108_0Output, mb_D_FF108_132MultiplierStage1Output);

    MB_D_FF_Float_108_132_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF108_132MultiplierStage1Output, mb_D_FF108_132MultiplierStage2Output);

    Multiplier_Float_108: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF108_132MultiplierStage2Output, flopocoMultiplier108WeightInput, Multiplier108_Output_132);

    MBRightSHR_Float_108_132: entity work.MBRightSHR(rtl)
    GENERIC MAP (43, NumberOfBits)
    PORT MAP (clk, rst, Multiplier108Weight, mbRightSHR108_132Output);

    MB_D_FF_Float_108_132_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR108_132Output, Multiplier108WeightOutput);

    InputIEEE_Float_108_132: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier108WeightOutput, flopocoMultiplier108WeightOutput);

    MB_D_FF_Float_108_132_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier108WeightOutput, flopocoMultiplier108WeightInput);

    MBRightSHR_Float_109_Input1133: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits)
    PORT MAP (clk, rst, Multiplier109Weight, mbRightSHR109_Input1_133Output);

    MB_D_FF_Float_109_133_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR109_Input1_133Output, Multiplier109WeightOutput);

    InputIEEE_Float_109_133: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier109WeightOutput, flopocoMultiplier109WeightOutput);

    MB_D_FF_Float_109_133_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier109WeightOutput, flopocoMultiplier109WeightInput);

    Multiplier_Float_109: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier109WeightInput, mb_D_FF109_133MultiplierStage2Output, Multiplier109_Output_133);

    MBRightSHR_Float_109_Input2_133: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR109_Input2_133Input, mbRightSHR109_Input2_133Output);

    MB_D_FF_Float_109_133_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR109_Input2_133Output, mb_D_FF109_133MultiplierStage1Output);

    MB_D_FF_Float_109_133_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF109_133MultiplierStage1Output, mb_D_FF109_133MultiplierStage2Output);

    MBRightSHR_Float_110_Input1134: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits)
    PORT MAP (clk, rst, Multiplier110Weight, mbRightSHR110_Input1_134Output);

    MB_D_FF_Float_110_134_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR110_Input1_134Output, Multiplier110WeightOutput);

    InputIEEE_Float_110_134: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier110WeightOutput, flopocoMultiplier110WeightOutput);

    MB_D_FF_Float_110_134_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier110WeightOutput, flopocoMultiplier110WeightInput);

    Multiplier_Float_110: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier110WeightInput, mb_D_FF110_134MultiplierStage2Output, Multiplier110_Output_134);

    MBRightSHR_Float_110_Input2_134: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR110_Input2_134Input, mbRightSHR110_Input2_134Output);

    MB_D_FF_Float_110_134_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR110_Input2_134Output, mb_D_FF110_134MultiplierStage1Output);

    MB_D_FF_Float_110_134_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF110_134MultiplierStage1Output, mb_D_FF110_134MultiplierStage2Output);

    MB_D_FF_Float_Adder18_Input1_24_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier110_Output_134, mb_D_FFAdder18_Input1_24_0Output);

    MB_D_FF_Float_24_135_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder18_Input1_24_0Output, mb_D_FF24_135AugendStage1Output);

    MB_D_FF_Float_24_135_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF24_135AugendStage1Output, mb_D_FF24_135AugendStage2Output);

    Adder_Float_24: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF24_135AugendStage2Output, mb_D_FF24_135AddendStage2Output, Adder24_Output_135);

    MB_D_FF_Float_Adder18_Input2_24_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier109_Output_133, mb_D_FFAdder18_Input2_24_0Output);

    MB_D_FF_Float_24_135_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder18_Input2_24_0Output, mb_D_FF24_135AddendStage1Output);

    MB_D_FF_Float_24_135_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF24_135AddendStage1Output, mb_D_FF24_135AddendStage2Output);

    MB_D_FF_Float_Multiplier17_Input1_111_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder24_Output_135, mb_D_FFMultiplier17_Input1_111_0Output);

    MB_D_FF_Float_111_136_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier17_Input1_111_0Output, mb_D_FF111_136MultiplicandStage1Output);

    MB_D_FF_Float_111_136_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF111_136MultiplicandStage1Output, mb_D_FF111_136MultiplicandStage2Output);

    Multiplier_Float_111: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF111_136MultiplicandStage2Output, mb_D_FF111_136MultiplierStage2Output, Multiplier111_Output_136);

    MB_D_FF_Float_Multiplier17_Input2_111_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier108_Output_132, mb_D_FFMultiplier17_Input2_111_0Output);

    MB_D_FF_Float_111_136_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier17_Input2_111_0Output, mb_D_FF111_136MultiplierStage1Output);

    MB_D_FF_Float_111_136_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF111_136MultiplierStage1Output, mb_D_FF111_136MultiplierStage2Output);

    MBRightSHR_Float_112_137: entity work.MBRightSHR(rtl)
    GENERIC MAP (4, NumberOfBits)
    PORT MAP (clk, rst, Multiplier112Weight, mbRightSHR112_137Output);

    MB_D_FF_Float_112_137_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR112_137Output, Multiplier112WeightOutput);

    InputIEEE_Float_112_137: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier112WeightOutput, flopocoMultiplier112WeightOutput);

    MB_D_FF_Float_112_137_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier112WeightOutput, flopocoMultiplier112WeightInput);

    Multiplier_Float_112: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier112WeightInput, mb_D_FF112_137MultiplierStage2Output, Multiplier112_Output_137);

    MB_D_FF_Float_Multiplier21_112_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier21_112_0Input, mb_D_FFMultiplier21_112_0Output);

    MB_D_FF_Float_112_137_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier21_112_0Output, mb_D_FF112_137MultiplierStage1Output);

    MB_D_FF_Float_112_137_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF112_137MultiplierStage1Output, mb_D_FF112_137MultiplierStage2Output);

    MBRightSHR_Float_113_138: entity work.MBRightSHR(rtl)
    GENERIC MAP (4, NumberOfBits)
    PORT MAP (clk, rst, Multiplier113Weight, mbRightSHR113_138Output);

    MB_D_FF_Float_113_138_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR113_138Output, Multiplier113WeightOutput);

    InputIEEE_Float_113_138: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier113WeightOutput, flopocoMultiplier113WeightOutput);

    MB_D_FF_Float_113_138_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier113WeightOutput, flopocoMultiplier113WeightInput);

    Multiplier_Float_113: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier113WeightInput, mb_D_FF113_138MultiplierStage2Output, Multiplier113_Output_138);

    MB_D_FF_Float_Multiplier21_113_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier21_113_0Input, mb_D_FFMultiplier21_113_0Output);

    MB_D_FF_Float_113_138_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier21_113_0Output, mb_D_FF113_138MultiplierStage1Output);

    MB_D_FF_Float_113_138_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF113_138MultiplierStage1Output, mb_D_FF113_138MultiplierStage2Output);

    MB_D_FF_Float_Adder20_Input1_25_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier113_Output_138, mb_D_FFAdder20_Input1_25_0Output);

    MB_D_FF_Float_25_139_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder20_Input1_25_0Output, mb_D_FF25_139AugendStage1Output);

    MB_D_FF_Float_25_139_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF25_139AugendStage1Output, mb_D_FF25_139AugendStage2Output);

    Adder_Float_25: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF25_139AugendStage2Output, mb_D_FF25_139AddendStage2Output, Adder25_Output_139);

    MB_D_FF_Float_Adder20_Input2_25_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier112_Output_137, mb_D_FFAdder20_Input2_25_0Output);

    MB_D_FF_Float_25_139_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder20_Input2_25_0Output, mb_D_FF25_139AddendStage1Output);

    MB_D_FF_Float_25_139_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF25_139AddendStage1Output, mb_D_FF25_139AddendStage2Output);

    MB_D_FF_Float_Multiplier19_114_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder25_Output_139, mb_D_FFMultiplier19_114_0Output);

    MB_D_FF_Float_114_140_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier19_114_0Output, mb_D_FF114_140MultiplierStage1Output);

    MB_D_FF_Float_114_140_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF114_140MultiplierStage1Output, mb_D_FF114_140MultiplierStage2Output);

    Multiplier_Float_114: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF114_140MultiplierStage2Output, mb_D_FF114_140MultiplicandStage2Output, Multiplier114_Output_140);

    MBRightSHR_Float_114_140: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR114_140Input, mbRightSHR114_140Output);

    MB_D_FF_Float_114_140_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR114_140Output, mb_D_FF114_140MultiplicandStage1Output);

    MB_D_FF_Float_114_140_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF114_140MultiplicandStage1Output, mb_D_FF114_140MultiplicandStage2Output);

    MB_D_FF_Float_Multiplier18_115_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier114_Output_140, mb_D_FFMultiplier18_115_0Output);

    MB_D_FF_Float_115_141_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier18_115_0Output, mb_D_FF115_141MultiplierStage1Output);

    MB_D_FF_Float_115_141_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF115_141MultiplierStage1Output, mb_D_FF115_141MultiplierStage2Output);

    Multiplier_Float_115: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF115_141MultiplierStage2Output, flopocoMultiplier115WeightInput, Multiplier115_Output_141);

    MBRightSHR_Float_115_141: entity work.MBRightSHR(rtl)
    GENERIC MAP (43, NumberOfBits)
    PORT MAP (clk, rst, Multiplier115Weight, mbRightSHR115_141Output);

    MB_D_FF_Float_115_141_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR115_141Output, Multiplier115WeightOutput);

    InputIEEE_Float_115_141: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier115WeightOutput, flopocoMultiplier115WeightOutput);

    MB_D_FF_Float_115_141_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier115WeightOutput, flopocoMultiplier115WeightInput);

    MBRightSHR_Float_116_Input1142: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits)
    PORT MAP (clk, rst, Multiplier116Weight, mbRightSHR116_Input1_142Output);

    MB_D_FF_Float_116_142_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR116_Input1_142Output, Multiplier116WeightOutput);

    InputIEEE_Float_116_142: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier116WeightOutput, flopocoMultiplier116WeightOutput);

    MB_D_FF_Float_116_142_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier116WeightOutput, flopocoMultiplier116WeightInput);

    Multiplier_Float_116: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier116WeightInput, mb_D_FF116_142MultiplierStage2Output, Multiplier116_Output_142);

    MBRightSHR_Float_116_Input2_142: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR116_Input2_142Input, mbRightSHR116_Input2_142Output);

    MB_D_FF_Float_116_142_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR116_Input2_142Output, mb_D_FF116_142MultiplierStage1Output);

    MB_D_FF_Float_116_142_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF116_142MultiplierStage1Output, mb_D_FF116_142MultiplierStage2Output);

    MBRightSHR_Float_117_Input1143: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits)
    PORT MAP (clk, rst, Multiplier117Weight, mbRightSHR117_Input1_143Output);

    MB_D_FF_Float_117_143_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR117_Input1_143Output, Multiplier117WeightOutput);

    InputIEEE_Float_117_143: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier117WeightOutput, flopocoMultiplier117WeightOutput);

    MB_D_FF_Float_117_143_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier117WeightOutput, flopocoMultiplier117WeightInput);

    Multiplier_Float_117: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier117WeightInput, mb_D_FF117_143MultiplierStage2Output, Multiplier117_Output_143);

    MBRightSHR_Float_117_Input2_143: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR117_Input2_143Input, mbRightSHR117_Input2_143Output);

    MB_D_FF_Float_117_143_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR117_Input2_143Output, mb_D_FF117_143MultiplierStage1Output);

    MB_D_FF_Float_117_143_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF117_143MultiplierStage1Output, mb_D_FF117_143MultiplierStage2Output);

    MB_D_FF_Float_Adder18_Input1_26_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier117_Output_143, mb_D_FFAdder18_Input1_26_0Output);

    MB_D_FF_Float_26_144_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder18_Input1_26_0Output, mb_D_FF26_144AugendStage1Output);

    MB_D_FF_Float_26_144_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF26_144AugendStage1Output, mb_D_FF26_144AugendStage2Output);

    Adder_Float_26: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF26_144AugendStage2Output, mb_D_FF26_144AddendStage2Output, Adder26_Output_144);

    MB_D_FF_Float_Adder18_Input2_26_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier116_Output_142, mb_D_FFAdder18_Input2_26_0Output);

    MB_D_FF_Float_26_144_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder18_Input2_26_0Output, mb_D_FF26_144AddendStage1Output);

    MB_D_FF_Float_26_144_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF26_144AddendStage1Output, mb_D_FF26_144AddendStage2Output);

    MB_D_FF_Float_Multiplier17_Input1_118_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder26_Output_144, mb_D_FFMultiplier17_Input1_118_0Output);

    MB_D_FF_Float_118_145_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier17_Input1_118_0Output, mb_D_FF118_145MultiplicandStage1Output);

    MB_D_FF_Float_118_145_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF118_145MultiplicandStage1Output, mb_D_FF118_145MultiplicandStage2Output);

    Multiplier_Float_118: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF118_145MultiplicandStage2Output, mb_D_FF118_145MultiplierStage2Output, Multiplier118_Output_145);

    MB_D_FF_Float_Multiplier17_Input2_118_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier115_Output_141, mb_D_FFMultiplier17_Input2_118_0Output);

    MB_D_FF_Float_118_145_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier17_Input2_118_0Output, mb_D_FF118_145MultiplierStage1Output);

    MB_D_FF_Float_118_145_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF118_145MultiplierStage1Output, mb_D_FF118_145MultiplierStage2Output);

    MB_D_FF_Float_Adder16_Input1_27_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier118_Output_145, mb_D_FFAdder16_Input1_27_0Output);

    MB_D_FF_Float_27_146_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder16_Input1_27_0Output, mb_D_FF27_146AugendStage1Output);

    MB_D_FF_Float_27_146_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF27_146AugendStage1Output, mb_D_FF27_146AugendStage2Output);

    Adder_Float_27: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF27_146AugendStage2Output, mb_D_FF27_146AddendStage2Output, Adder27_Output_146);

    MB_D_FF_Float_Adder16_Input2_27_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier111_Output_136, mb_D_FFAdder16_Input2_27_0Output);

    MB_D_FF_Float_27_146_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder16_Input2_27_0Output, mb_D_FF27_146AddendStage1Output);

    MB_D_FF_Float_27_146_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF27_146AddendStage1Output, mb_D_FF27_146AddendStage2Output);

    MB_D_FF_Float_Multiplier15_119_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder27_Output_146, mb_D_FFMultiplier15_119_0Output);

    MB_D_FF_Float_119_147_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier15_119_0Output, mb_D_FF119_147MultiplierStage1Output);

    MB_D_FF_Float_119_147_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF119_147MultiplierStage1Output, mb_D_FF119_147MultiplierStage2Output);

    Multiplier_Float_119: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF119_147MultiplierStage2Output, mb_D_FF119_147MultiplicandStage2Output, Multiplier119_Output_147);

    MBRightSHR_Float_119_147: entity work.MBRightSHR(rtl)
    GENERIC MAP (82, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR119_147Input, mbRightSHR119_147Output);

    MB_D_FF_Float_119_147_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR119_147Output, mb_D_FF119_147MultiplicandStage1Output);

    MB_D_FF_Float_119_147_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF119_147MultiplicandStage1Output, mb_D_FF119_147MultiplicandStage2Output);

    MB_D_FF_Float_Multiplier14_120_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier119_Output_147, mb_D_FFMultiplier14_120_0Output);

    MB_D_FF_Float_120_148_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier14_120_0Output, mb_D_FF120_148MultiplierStage1Output);

    MB_D_FF_Float_120_148_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF120_148MultiplierStage1Output, mb_D_FF120_148MultiplierStage2Output);

    Multiplier_Float_120: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF120_148MultiplierStage2Output, flopocoMultiplier120WeightInput, Multiplier120_Output_148);

    MBRightSHR_Float_120_148: entity work.MBRightSHR(rtl)
    GENERIC MAP (89, NumberOfBits)
    PORT MAP (clk, rst, Multiplier120Weight, mbRightSHR120_148Output);

    MB_D_FF_Float_120_148_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR120_148Output, Multiplier120WeightOutput);

    InputIEEE_Float_120_148: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier120WeightOutput, flopocoMultiplier120WeightOutput);

    MB_D_FF_Float_120_148_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier120WeightOutput, flopocoMultiplier120WeightInput);

    MBRightSHR_Float_121_149: entity work.MBRightSHR(rtl)
    GENERIC MAP (4, NumberOfBits)
    PORT MAP (clk, rst, Multiplier121Weight, mbRightSHR121_149Output);

    MB_D_FF_Float_121_149_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR121_149Output, Multiplier121WeightOutput);

    InputIEEE_Float_121_149: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier121WeightOutput, flopocoMultiplier121WeightOutput);

    MB_D_FF_Float_121_149_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier121WeightOutput, flopocoMultiplier121WeightInput);

    Multiplier_Float_121: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier121WeightInput, mb_D_FF121_149MultiplierStage2Output, Multiplier121_Output_149);

    MB_D_FF_Float_Multiplier21_121_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier21_121_0Input, mb_D_FFMultiplier21_121_0Output);

    MB_D_FF_Float_121_149_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier21_121_0Output, mb_D_FF121_149MultiplierStage1Output);

    MB_D_FF_Float_121_149_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF121_149MultiplierStage1Output, mb_D_FF121_149MultiplierStage2Output);

    MBRightSHR_Float_122_150: entity work.MBRightSHR(rtl)
    GENERIC MAP (4, NumberOfBits)
    PORT MAP (clk, rst, Multiplier122Weight, mbRightSHR122_150Output);

    MB_D_FF_Float_122_150_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR122_150Output, Multiplier122WeightOutput);

    InputIEEE_Float_122_150: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier122WeightOutput, flopocoMultiplier122WeightOutput);

    MB_D_FF_Float_122_150_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier122WeightOutput, flopocoMultiplier122WeightInput);

    Multiplier_Float_122: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier122WeightInput, mb_D_FF122_150MultiplierStage2Output, Multiplier122_Output_150);

    MB_D_FF_Float_Multiplier21_122_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier21_122_0Input, mb_D_FFMultiplier21_122_0Output);

    MB_D_FF_Float_122_150_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier21_122_0Output, mb_D_FF122_150MultiplierStage1Output);

    MB_D_FF_Float_122_150_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF122_150MultiplierStage1Output, mb_D_FF122_150MultiplierStage2Output);

    MB_D_FF_Float_Adder20_Input1_28_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier122_Output_150, mb_D_FFAdder20_Input1_28_0Output);

    MB_D_FF_Float_28_151_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder20_Input1_28_0Output, mb_D_FF28_151AugendStage1Output);

    MB_D_FF_Float_28_151_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF28_151AugendStage1Output, mb_D_FF28_151AugendStage2Output);

    Adder_Float_28: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF28_151AugendStage2Output, mb_D_FF28_151AddendStage2Output, Adder28_Output_151);

    MB_D_FF_Float_Adder20_Input2_28_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier121_Output_149, mb_D_FFAdder20_Input2_28_0Output);

    MB_D_FF_Float_28_151_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder20_Input2_28_0Output, mb_D_FF28_151AddendStage1Output);

    MB_D_FF_Float_28_151_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF28_151AddendStage1Output, mb_D_FF28_151AddendStage2Output);

    MB_D_FF_Float_Multiplier19_123_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder28_Output_151, mb_D_FFMultiplier19_123_0Output);

    MB_D_FF_Float_123_152_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier19_123_0Output, mb_D_FF123_152MultiplierStage1Output);

    MB_D_FF_Float_123_152_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF123_152MultiplierStage1Output, mb_D_FF123_152MultiplierStage2Output);

    Multiplier_Float_123: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF123_152MultiplierStage2Output, mb_D_FF123_152MultiplicandStage2Output, Multiplier123_Output_152);

    MBRightSHR_Float_123_152: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR123_152Input, mbRightSHR123_152Output);

    MB_D_FF_Float_123_152_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR123_152Output, mb_D_FF123_152MultiplicandStage1Output);

    MB_D_FF_Float_123_152_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF123_152MultiplicandStage1Output, mb_D_FF123_152MultiplicandStage2Output);

    MB_D_FF_Float_Multiplier18_124_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier123_Output_152, mb_D_FFMultiplier18_124_0Output);

    MB_D_FF_Float_124_153_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier18_124_0Output, mb_D_FF124_153MultiplierStage1Output);

    MB_D_FF_Float_124_153_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF124_153MultiplierStage1Output, mb_D_FF124_153MultiplierStage2Output);

    Multiplier_Float_124: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF124_153MultiplierStage2Output, flopocoMultiplier124WeightInput, Multiplier124_Output_153);

    MBRightSHR_Float_124_153: entity work.MBRightSHR(rtl)
    GENERIC MAP (43, NumberOfBits)
    PORT MAP (clk, rst, Multiplier124Weight, mbRightSHR124_153Output);

    MB_D_FF_Float_124_153_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR124_153Output, Multiplier124WeightOutput);

    InputIEEE_Float_124_153: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier124WeightOutput, flopocoMultiplier124WeightOutput);

    MB_D_FF_Float_124_153_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier124WeightOutput, flopocoMultiplier124WeightInput);

    MBRightSHR_Float_125_Input1154: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits)
    PORT MAP (clk, rst, Multiplier125Weight, mbRightSHR125_Input1_154Output);

    MB_D_FF_Float_125_154_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR125_Input1_154Output, Multiplier125WeightOutput);

    InputIEEE_Float_125_154: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier125WeightOutput, flopocoMultiplier125WeightOutput);

    MB_D_FF_Float_125_154_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier125WeightOutput, flopocoMultiplier125WeightInput);

    Multiplier_Float_125: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier125WeightInput, mb_D_FF125_154MultiplierStage2Output, Multiplier125_Output_154);

    MBRightSHR_Float_125_Input2_154: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR125_Input2_154Input, mbRightSHR125_Input2_154Output);

    MB_D_FF_Float_125_154_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR125_Input2_154Output, mb_D_FF125_154MultiplierStage1Output);

    MB_D_FF_Float_125_154_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF125_154MultiplierStage1Output, mb_D_FF125_154MultiplierStage2Output);

    MBRightSHR_Float_126_Input1155: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits)
    PORT MAP (clk, rst, Multiplier126Weight, mbRightSHR126_Input1_155Output);

    MB_D_FF_Float_126_155_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR126_Input1_155Output, Multiplier126WeightOutput);

    InputIEEE_Float_126_155: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier126WeightOutput, flopocoMultiplier126WeightOutput);

    MB_D_FF_Float_126_155_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier126WeightOutput, flopocoMultiplier126WeightInput);

    Multiplier_Float_126: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier126WeightInput, mb_D_FF126_155MultiplierStage2Output, Multiplier126_Output_155);

    MBRightSHR_Float_126_Input2_155: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR126_Input2_155Input, mbRightSHR126_Input2_155Output);

    MB_D_FF_Float_126_155_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR126_Input2_155Output, mb_D_FF126_155MultiplierStage1Output);

    MB_D_FF_Float_126_155_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF126_155MultiplierStage1Output, mb_D_FF126_155MultiplierStage2Output);

    MB_D_FF_Float_Adder18_Input1_29_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier126_Output_155, mb_D_FFAdder18_Input1_29_0Output);

    MB_D_FF_Float_29_156_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder18_Input1_29_0Output, mb_D_FF29_156AugendStage1Output);

    MB_D_FF_Float_29_156_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF29_156AugendStage1Output, mb_D_FF29_156AugendStage2Output);

    Adder_Float_29: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF29_156AugendStage2Output, mb_D_FF29_156AddendStage2Output, Adder29_Output_156);

    MB_D_FF_Float_Adder18_Input2_29_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier125_Output_154, mb_D_FFAdder18_Input2_29_0Output);

    MB_D_FF_Float_29_156_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder18_Input2_29_0Output, mb_D_FF29_156AddendStage1Output);

    MB_D_FF_Float_29_156_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF29_156AddendStage1Output, mb_D_FF29_156AddendStage2Output);

    MB_D_FF_Float_Multiplier17_Input1_127_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder29_Output_156, mb_D_FFMultiplier17_Input1_127_0Output);

    MB_D_FF_Float_127_157_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier17_Input1_127_0Output, mb_D_FF127_157MultiplicandStage1Output);

    MB_D_FF_Float_127_157_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF127_157MultiplicandStage1Output, mb_D_FF127_157MultiplicandStage2Output);

    Multiplier_Float_127: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF127_157MultiplicandStage2Output, mb_D_FF127_157MultiplierStage2Output, Multiplier127_Output_157);

    MB_D_FF_Float_Multiplier17_Input2_127_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier124_Output_153, mb_D_FFMultiplier17_Input2_127_0Output);

    MB_D_FF_Float_127_157_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier17_Input2_127_0Output, mb_D_FF127_157MultiplierStage1Output);

    MB_D_FF_Float_127_157_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF127_157MultiplierStage1Output, mb_D_FF127_157MultiplierStage2Output);

    MBRightSHR_Float_128_158: entity work.MBRightSHR(rtl)
    GENERIC MAP (4, NumberOfBits)
    PORT MAP (clk, rst, Multiplier128Weight, mbRightSHR128_158Output);

    MB_D_FF_Float_128_158_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR128_158Output, Multiplier128WeightOutput);

    InputIEEE_Float_128_158: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier128WeightOutput, flopocoMultiplier128WeightOutput);

    MB_D_FF_Float_128_158_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier128WeightOutput, flopocoMultiplier128WeightInput);

    Multiplier_Float_128: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier128WeightInput, mb_D_FF128_158MultiplierStage2Output, Multiplier128_Output_158);

    MB_D_FF_Float_Multiplier21_128_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier21_128_0Input, mb_D_FFMultiplier21_128_0Output);

    MB_D_FF_Float_128_158_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier21_128_0Output, mb_D_FF128_158MultiplierStage1Output);

    MB_D_FF_Float_128_158_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF128_158MultiplierStage1Output, mb_D_FF128_158MultiplierStage2Output);

    MBRightSHR_Float_129_159: entity work.MBRightSHR(rtl)
    GENERIC MAP (4, NumberOfBits)
    PORT MAP (clk, rst, Multiplier129Weight, mbRightSHR129_159Output);

    MB_D_FF_Float_129_159_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR129_159Output, Multiplier129WeightOutput);

    InputIEEE_Float_129_159: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier129WeightOutput, flopocoMultiplier129WeightOutput);

    MB_D_FF_Float_129_159_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier129WeightOutput, flopocoMultiplier129WeightInput);

    Multiplier_Float_129: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier129WeightInput, mb_D_FF129_159MultiplierStage2Output, Multiplier129_Output_159);

    MB_D_FF_Float_Multiplier21_129_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier21_129_0Input, mb_D_FFMultiplier21_129_0Output);

    MB_D_FF_Float_129_159_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier21_129_0Output, mb_D_FF129_159MultiplierStage1Output);

    MB_D_FF_Float_129_159_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF129_159MultiplierStage1Output, mb_D_FF129_159MultiplierStage2Output);

    MB_D_FF_Float_Adder20_Input1_30_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier129_Output_159, mb_D_FFAdder20_Input1_30_0Output);

    MB_D_FF_Float_30_160_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder20_Input1_30_0Output, mb_D_FF30_160AugendStage1Output);

    MB_D_FF_Float_30_160_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF30_160AugendStage1Output, mb_D_FF30_160AugendStage2Output);

    Adder_Float_30: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF30_160AugendStage2Output, mb_D_FF30_160AddendStage2Output, Adder30_Output_160);

    MB_D_FF_Float_Adder20_Input2_30_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier128_Output_158, mb_D_FFAdder20_Input2_30_0Output);

    MB_D_FF_Float_30_160_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder20_Input2_30_0Output, mb_D_FF30_160AddendStage1Output);

    MB_D_FF_Float_30_160_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF30_160AddendStage1Output, mb_D_FF30_160AddendStage2Output);

    MB_D_FF_Float_Multiplier19_130_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder30_Output_160, mb_D_FFMultiplier19_130_0Output);

    MB_D_FF_Float_130_161_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier19_130_0Output, mb_D_FF130_161MultiplierStage1Output);

    MB_D_FF_Float_130_161_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF130_161MultiplierStage1Output, mb_D_FF130_161MultiplierStage2Output);

    Multiplier_Float_130: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF130_161MultiplierStage2Output, mb_D_FF130_161MultiplicandStage2Output, Multiplier130_Output_161);

    MBRightSHR_Float_130_161: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR130_161Input, mbRightSHR130_161Output);

    MB_D_FF_Float_130_161_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR130_161Output, mb_D_FF130_161MultiplicandStage1Output);

    MB_D_FF_Float_130_161_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF130_161MultiplicandStage1Output, mb_D_FF130_161MultiplicandStage2Output);

    MB_D_FF_Float_Multiplier18_131_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier130_Output_161, mb_D_FFMultiplier18_131_0Output);

    MB_D_FF_Float_131_162_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier18_131_0Output, mb_D_FF131_162MultiplierStage1Output);

    MB_D_FF_Float_131_162_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF131_162MultiplierStage1Output, mb_D_FF131_162MultiplierStage2Output);

    Multiplier_Float_131: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF131_162MultiplierStage2Output, flopocoMultiplier131WeightInput, Multiplier131_Output_162);

    MBRightSHR_Float_131_162: entity work.MBRightSHR(rtl)
    GENERIC MAP (43, NumberOfBits)
    PORT MAP (clk, rst, Multiplier131Weight, mbRightSHR131_162Output);

    MB_D_FF_Float_131_162_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR131_162Output, Multiplier131WeightOutput);

    InputIEEE_Float_131_162: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier131WeightOutput, flopocoMultiplier131WeightOutput);

    MB_D_FF_Float_131_162_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier131WeightOutput, flopocoMultiplier131WeightInput);

    MBRightSHR_Float_132_Input1163: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits)
    PORT MAP (clk, rst, Multiplier132Weight, mbRightSHR132_Input1_163Output);

    MB_D_FF_Float_132_163_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR132_Input1_163Output, Multiplier132WeightOutput);

    InputIEEE_Float_132_163: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier132WeightOutput, flopocoMultiplier132WeightOutput);

    MB_D_FF_Float_132_163_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier132WeightOutput, flopocoMultiplier132WeightInput);

    Multiplier_Float_132: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier132WeightInput, mb_D_FF132_163MultiplierStage2Output, Multiplier132_Output_163);

    MBRightSHR_Float_132_Input2_163: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR132_Input2_163Input, mbRightSHR132_Input2_163Output);

    MB_D_FF_Float_132_163_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR132_Input2_163Output, mb_D_FF132_163MultiplierStage1Output);

    MB_D_FF_Float_132_163_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF132_163MultiplierStage1Output, mb_D_FF132_163MultiplierStage2Output);

    MBRightSHR_Float_133_Input1164: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits)
    PORT MAP (clk, rst, Multiplier133Weight, mbRightSHR133_Input1_164Output);

    MB_D_FF_Float_133_164_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR133_Input1_164Output, Multiplier133WeightOutput);

    InputIEEE_Float_133_164: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier133WeightOutput, flopocoMultiplier133WeightOutput);

    MB_D_FF_Float_133_164_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier133WeightOutput, flopocoMultiplier133WeightInput);

    Multiplier_Float_133: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier133WeightInput, mb_D_FF133_164MultiplierStage2Output, Multiplier133_Output_164);

    MBRightSHR_Float_133_Input2_164: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR133_Input2_164Input, mbRightSHR133_Input2_164Output);

    MB_D_FF_Float_133_164_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR133_Input2_164Output, mb_D_FF133_164MultiplierStage1Output);

    MB_D_FF_Float_133_164_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF133_164MultiplierStage1Output, mb_D_FF133_164MultiplierStage2Output);

    MB_D_FF_Float_Adder18_Input1_31_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier133_Output_164, mb_D_FFAdder18_Input1_31_0Output);

    MB_D_FF_Float_31_165_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder18_Input1_31_0Output, mb_D_FF31_165AugendStage1Output);

    MB_D_FF_Float_31_165_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF31_165AugendStage1Output, mb_D_FF31_165AugendStage2Output);

    Adder_Float_31: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF31_165AugendStage2Output, mb_D_FF31_165AddendStage2Output, Adder31_Output_165);

    MB_D_FF_Float_Adder18_Input2_31_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier132_Output_163, mb_D_FFAdder18_Input2_31_0Output);

    MB_D_FF_Float_31_165_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder18_Input2_31_0Output, mb_D_FF31_165AddendStage1Output);

    MB_D_FF_Float_31_165_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF31_165AddendStage1Output, mb_D_FF31_165AddendStage2Output);

    MB_D_FF_Float_Multiplier17_Input1_134_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder31_Output_165, mb_D_FFMultiplier17_Input1_134_0Output);

    MB_D_FF_Float_134_166_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier17_Input1_134_0Output, mb_D_FF134_166MultiplicandStage1Output);

    MB_D_FF_Float_134_166_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF134_166MultiplicandStage1Output, mb_D_FF134_166MultiplicandStage2Output);

    Multiplier_Float_134: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF134_166MultiplicandStage2Output, mb_D_FF134_166MultiplierStage2Output, Multiplier134_Output_166);

    MB_D_FF_Float_Multiplier17_Input2_134_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier131_Output_162, mb_D_FFMultiplier17_Input2_134_0Output);

    MB_D_FF_Float_134_166_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier17_Input2_134_0Output, mb_D_FF134_166MultiplierStage1Output);

    MB_D_FF_Float_134_166_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF134_166MultiplierStage1Output, mb_D_FF134_166MultiplierStage2Output);

    MB_D_FF_Float_Adder16_Input1_32_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier134_Output_166, mb_D_FFAdder16_Input1_32_0Output);

    MB_D_FF_Float_32_167_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder16_Input1_32_0Output, mb_D_FF32_167AugendStage1Output);

    MB_D_FF_Float_32_167_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF32_167AugendStage1Output, mb_D_FF32_167AugendStage2Output);

    Adder_Float_32: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF32_167AugendStage2Output, mb_D_FF32_167AddendStage2Output, Adder32_Output_167);

    MB_D_FF_Float_Adder16_Input2_32_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier127_Output_157, mb_D_FFAdder16_Input2_32_0Output);

    MB_D_FF_Float_32_167_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder16_Input2_32_0Output, mb_D_FF32_167AddendStage1Output);

    MB_D_FF_Float_32_167_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF32_167AddendStage1Output, mb_D_FF32_167AddendStage2Output);

    MB_D_FF_Float_Multiplier15_135_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder32_Output_167, mb_D_FFMultiplier15_135_0Output);

    MB_D_FF_Float_135_168_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier15_135_0Output, mb_D_FF135_168MultiplierStage1Output);

    MB_D_FF_Float_135_168_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF135_168MultiplierStage1Output, mb_D_FF135_168MultiplierStage2Output);

    Multiplier_Float_135: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF135_168MultiplierStage2Output, mb_D_FF135_168MultiplicandStage2Output, Multiplier135_Output_168);

    MBRightSHR_Float_135_168: entity work.MBRightSHR(rtl)
    GENERIC MAP (82, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR135_168Input, mbRightSHR135_168Output);

    MB_D_FF_Float_135_168_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR135_168Output, mb_D_FF135_168MultiplicandStage1Output);

    MB_D_FF_Float_135_168_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF135_168MultiplicandStage1Output, mb_D_FF135_168MultiplicandStage2Output);

    MB_D_FF_Float_Multiplier14_136_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier135_Output_168, mb_D_FFMultiplier14_136_0Output);

    MB_D_FF_Float_136_169_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier14_136_0Output, mb_D_FF136_169MultiplierStage1Output);

    MB_D_FF_Float_136_169_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF136_169MultiplierStage1Output, mb_D_FF136_169MultiplierStage2Output);

    Multiplier_Float_136: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF136_169MultiplierStage2Output, flopocoMultiplier136WeightInput, Multiplier136_Output_169);

    MBRightSHR_Float_136_169: entity work.MBRightSHR(rtl)
    GENERIC MAP (89, NumberOfBits)
    PORT MAP (clk, rst, Multiplier136Weight, mbRightSHR136_169Output);

    MB_D_FF_Float_136_169_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR136_169Output, Multiplier136WeightOutput);

    InputIEEE_Float_136_169: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier136WeightOutput, flopocoMultiplier136WeightOutput);

    MB_D_FF_Float_136_169_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier136WeightOutput, flopocoMultiplier136WeightInput);

    MB_D_FF_Float_Adder13_Input1_33_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier136_Output_169, mb_D_FFAdder13_Input1_33_0Output);

    MB_D_FF_Float_33_170_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder13_Input1_33_0Output, mb_D_FF33_170AugendStage1Output);

    MB_D_FF_Float_33_170_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF33_170AugendStage1Output, mb_D_FF33_170AugendStage2Output);

    Adder_Float_33: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF33_170AugendStage2Output, mb_D_FF33_170AddendStage2Output, Adder33_Output_170);

    MB_D_FF_Float_Adder13_Input2_33_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier120_Output_148, mb_D_FFAdder13_Input2_33_0Output);

    MB_D_FF_Float_33_170_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder13_Input2_33_0Output, mb_D_FF33_170AddendStage1Output);

    MB_D_FF_Float_33_170_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF33_170AddendStage1Output, mb_D_FF33_170AddendStage2Output);

    MB_D_FF_Float_Multiplier12_137_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder33_Output_170, mb_D_FFMultiplier12_137_0Output);

    MB_D_FF_Float_137_171_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier12_137_0Output, mb_D_FF137_171MultiplierStage1Output);

    MB_D_FF_Float_137_171_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF137_171MultiplierStage1Output, mb_D_FF137_171MultiplierStage2Output);

    Multiplier_Float_137: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF137_171MultiplierStage2Output, mb_D_FF137_171MultiplicandStage2Output, Multiplier137_Output_171);

    MBRightSHR_Float_137_171: entity work.MBRightSHR(rtl)
    GENERIC MAP (121, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR137_171Input, mbRightSHR137_171Output);

    MB_D_FF_Float_137_171_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR137_171Output, mb_D_FF137_171MultiplicandStage1Output);

    MB_D_FF_Float_137_171_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF137_171MultiplicandStage1Output, mb_D_FF137_171MultiplicandStage2Output);

    MBRightSHR_Float_138_Input1172: entity work.MBRightSHR(rtl)
    GENERIC MAP (50, NumberOfBits)
    PORT MAP (clk, rst, Multiplier138Weight, mbRightSHR138_Input1_172Output);

    MB_D_FF_Float_138_172_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR138_Input1_172Output, Multiplier138WeightOutput);

    InputIEEE_Float_138_172: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier138WeightOutput, flopocoMultiplier138WeightOutput);

    MB_D_FF_Float_138_172_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier138WeightOutput, flopocoMultiplier138WeightInput);

    Multiplier_Float_138: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier138WeightInput, mb_D_FF138_172MultiplierStage2Output, Multiplier138_Output_172);

    MBRightSHR_Float_138_Input2_172: entity work.MBRightSHR(rtl)
    GENERIC MAP (50, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR138_Input2_172Input, mbRightSHR138_Input2_172Output);

    MB_D_FF_Float_138_172_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR138_Input2_172Output, mb_D_FF138_172MultiplierStage1Output);

    MB_D_FF_Float_138_172_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF138_172MultiplierStage1Output, mb_D_FF138_172MultiplierStage2Output);

    MBRightSHR_Float_139_Input1173: entity work.MBRightSHR(rtl)
    GENERIC MAP (50, NumberOfBits)
    PORT MAP (clk, rst, Multiplier139Weight, mbRightSHR139_Input1_173Output);

    MB_D_FF_Float_139_173_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR139_Input1_173Output, Multiplier139WeightOutput);

    InputIEEE_Float_139_173: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier139WeightOutput, flopocoMultiplier139WeightOutput);

    MB_D_FF_Float_139_173_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier139WeightOutput, flopocoMultiplier139WeightInput);

    Multiplier_Float_139: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier139WeightInput, mb_D_FF139_173MultiplierStage2Output, Multiplier139_Output_173);

    MBRightSHR_Float_139_Input2_173: entity work.MBRightSHR(rtl)
    GENERIC MAP (50, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR139_Input2_173Input, mbRightSHR139_Input2_173Output);

    MB_D_FF_Float_139_173_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR139_Input2_173Output, mb_D_FF139_173MultiplierStage1Output);

    MB_D_FF_Float_139_173_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF139_173MultiplierStage1Output, mb_D_FF139_173MultiplierStage2Output);

    MB_D_FF_Float_Adder16_Input1_34_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier139_Output_173, mb_D_FFAdder16_Input1_34_0Output);

    MB_D_FF_Float_34_174_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder16_Input1_34_0Output, mb_D_FF34_174AugendStage1Output);

    MB_D_FF_Float_34_174_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF34_174AugendStage1Output, mb_D_FF34_174AugendStage2Output);

    Adder_Float_34: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF34_174AugendStage2Output, mb_D_FF34_174AddendStage2Output, Adder34_Output_174);

    MB_D_FF_Float_Adder16_Input2_34_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier138_Output_172, mb_D_FFAdder16_Input2_34_0Output);

    MB_D_FF_Float_34_174_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder16_Input2_34_0Output, mb_D_FF34_174AddendStage1Output);

    MB_D_FF_Float_34_174_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF34_174AddendStage1Output, mb_D_FF34_174AddendStage2Output);

    MB_D_FF_Float_Multiplier15_140_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder34_Output_174, mb_D_FFMultiplier15_140_0Output);

    MB_D_FF_Float_140_175_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier15_140_0Output, mb_D_FF140_175MultiplierStage1Output);

    MB_D_FF_Float_140_175_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF140_175MultiplierStage1Output, mb_D_FF140_175MultiplierStage2Output);

    Multiplier_Float_140: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF140_175MultiplierStage2Output, mb_D_FF140_175MultiplicandStage2Output, Multiplier140_Output_175);

    MBRightSHR_Float_140_175: entity work.MBRightSHR(rtl)
    GENERIC MAP (82, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR140_175Input, mbRightSHR140_175Output);

    MB_D_FF_Float_140_175_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR140_175Output, mb_D_FF140_175MultiplicandStage1Output);

    MB_D_FF_Float_140_175_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF140_175MultiplicandStage1Output, mb_D_FF140_175MultiplicandStage2Output);

    MB_D_FF_Float_Multiplier14_141_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier140_Output_175, mb_D_FFMultiplier14_141_0Output);

    MB_D_FF_Float_141_176_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier14_141_0Output, mb_D_FF141_176MultiplierStage1Output);

    MB_D_FF_Float_141_176_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF141_176MultiplierStage1Output, mb_D_FF141_176MultiplierStage2Output);

    Multiplier_Float_141: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF141_176MultiplierStage2Output, flopocoMultiplier141WeightInput, Multiplier141_Output_176);

    MBRightSHR_Float_141_176: entity work.MBRightSHR(rtl)
    GENERIC MAP (89, NumberOfBits)
    PORT MAP (clk, rst, Multiplier141Weight, mbRightSHR141_176Output);

    MB_D_FF_Float_141_176_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR141_176Output, Multiplier141WeightOutput);

    InputIEEE_Float_141_176: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier141WeightOutput, flopocoMultiplier141WeightOutput);

    MB_D_FF_Float_141_176_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier141WeightOutput, flopocoMultiplier141WeightInput);

    MB_D_FF_Float_Multiplier13_142_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier141_Output_176, mb_D_FFMultiplier13_142_0Output);

    MB_D_FF_Float_142_177_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier13_142_0Output, mb_D_FF142_177MultiplierStage1Output);

    MB_D_FF_Float_142_177_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF142_177MultiplierStage1Output, mb_D_FF142_177MultiplierStage2Output);

    Multiplier_Float_142: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF142_177MultiplierStage2Output, flopocoMultiplier142WeightInput, Multiplier142_Output_177);

    MBRightSHR_Float_142_177: entity work.MBRightSHR(rtl)
    GENERIC MAP (96, NumberOfBits)
    PORT MAP (clk, rst, Multiplier142Weight, mbRightSHR142_177Output);

    MB_D_FF_Float_142_177_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR142_177Output, Multiplier142WeightOutput);

    InputIEEE_Float_142_177: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier142WeightOutput, flopocoMultiplier142WeightOutput);

    MB_D_FF_Float_142_177_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier142WeightOutput, flopocoMultiplier142WeightInput);

    MBRightSHR_Float_143_Input1178: entity work.MBRightSHR(rtl)
    GENERIC MAP (50, NumberOfBits)
    PORT MAP (clk, rst, Multiplier143Weight, mbRightSHR143_Input1_178Output);

    MB_D_FF_Float_143_178_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR143_Input1_178Output, Multiplier143WeightOutput);

    InputIEEE_Float_143_178: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier143WeightOutput, flopocoMultiplier143WeightOutput);

    MB_D_FF_Float_143_178_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier143WeightOutput, flopocoMultiplier143WeightInput);

    Multiplier_Float_143: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier143WeightInput, mb_D_FF143_178MultiplierStage2Output, Multiplier143_Output_178);

    MBRightSHR_Float_143_Input2_178: entity work.MBRightSHR(rtl)
    GENERIC MAP (50, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR143_Input2_178Input, mbRightSHR143_Input2_178Output);

    MB_D_FF_Float_143_178_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR143_Input2_178Output, mb_D_FF143_178MultiplierStage1Output);

    MB_D_FF_Float_143_178_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF143_178MultiplierStage1Output, mb_D_FF143_178MultiplierStage2Output);

    MBRightSHR_Float_144_Input1179: entity work.MBRightSHR(rtl)
    GENERIC MAP (50, NumberOfBits)
    PORT MAP (clk, rst, Multiplier144Weight, mbRightSHR144_Input1_179Output);

    MB_D_FF_Float_144_179_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR144_Input1_179Output, Multiplier144WeightOutput);

    InputIEEE_Float_144_179: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier144WeightOutput, flopocoMultiplier144WeightOutput);

    MB_D_FF_Float_144_179_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier144WeightOutput, flopocoMultiplier144WeightInput);

    Multiplier_Float_144: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier144WeightInput, mb_D_FF144_179MultiplierStage2Output, Multiplier144_Output_179);

    MBRightSHR_Float_144_Input2_179: entity work.MBRightSHR(rtl)
    GENERIC MAP (50, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR144_Input2_179Input, mbRightSHR144_Input2_179Output);

    MB_D_FF_Float_144_179_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR144_Input2_179Output, mb_D_FF144_179MultiplierStage1Output);

    MB_D_FF_Float_144_179_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF144_179MultiplierStage1Output, mb_D_FF144_179MultiplierStage2Output);

    MB_D_FF_Float_Adder16_Input1_35_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier144_Output_179, mb_D_FFAdder16_Input1_35_0Output);

    MB_D_FF_Float_35_180_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder16_Input1_35_0Output, mb_D_FF35_180AugendStage1Output);

    MB_D_FF_Float_35_180_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF35_180AugendStage1Output, mb_D_FF35_180AugendStage2Output);

    Adder_Float_35: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF35_180AugendStage2Output, mb_D_FF35_180AddendStage2Output, Adder35_Output_180);

    MB_D_FF_Float_Adder16_Input2_35_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier143_Output_178, mb_D_FFAdder16_Input2_35_0Output);

    MB_D_FF_Float_35_180_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder16_Input2_35_0Output, mb_D_FF35_180AddendStage1Output);

    MB_D_FF_Float_35_180_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF35_180AddendStage1Output, mb_D_FF35_180AddendStage2Output);

    MB_D_FF_Float_Multiplier15_145_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder35_Output_180, mb_D_FFMultiplier15_145_0Output);

    MB_D_FF_Float_145_181_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier15_145_0Output, mb_D_FF145_181MultiplierStage1Output);

    MB_D_FF_Float_145_181_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF145_181MultiplierStage1Output, mb_D_FF145_181MultiplierStage2Output);

    Multiplier_Float_145: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF145_181MultiplierStage2Output, mb_D_FF145_181MultiplicandStage2Output, Multiplier145_Output_181);

    MBRightSHR_Float_145_181: entity work.MBRightSHR(rtl)
    GENERIC MAP (82, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR145_181Input, mbRightSHR145_181Output);

    MB_D_FF_Float_145_181_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR145_181Output, mb_D_FF145_181MultiplicandStage1Output);

    MB_D_FF_Float_145_181_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF145_181MultiplicandStage1Output, mb_D_FF145_181MultiplicandStage2Output);

    MB_D_FF_Float_Multiplier14_146_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier145_Output_181, mb_D_FFMultiplier14_146_0Output);

    MB_D_FF_Float_146_182_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier14_146_0Output, mb_D_FF146_182MultiplierStage1Output);

    MB_D_FF_Float_146_182_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF146_182MultiplierStage1Output, mb_D_FF146_182MultiplierStage2Output);

    Multiplier_Float_146: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF146_182MultiplierStage2Output, flopocoMultiplier146WeightInput, Multiplier146_Output_182);

    MBRightSHR_Float_146_182: entity work.MBRightSHR(rtl)
    GENERIC MAP (89, NumberOfBits)
    PORT MAP (clk, rst, Multiplier146Weight, mbRightSHR146_182Output);

    MB_D_FF_Float_146_182_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR146_182Output, Multiplier146WeightOutput);

    InputIEEE_Float_146_182: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier146WeightOutput, flopocoMultiplier146WeightOutput);

    MB_D_FF_Float_146_182_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier146WeightOutput, flopocoMultiplier146WeightInput);

    MB_D_FF_Float_Multiplier13_147_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier146_Output_182, mb_D_FFMultiplier13_147_0Output);

    MB_D_FF_Float_147_183_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier13_147_0Output, mb_D_FF147_183MultiplierStage1Output);

    MB_D_FF_Float_147_183_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF147_183MultiplierStage1Output, mb_D_FF147_183MultiplierStage2Output);

    Multiplier_Float_147: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF147_183MultiplierStage2Output, flopocoMultiplier147WeightInput, Multiplier147_Output_183);

    MBRightSHR_Float_147_183: entity work.MBRightSHR(rtl)
    GENERIC MAP (96, NumberOfBits)
    PORT MAP (clk, rst, Multiplier147Weight, mbRightSHR147_183Output);

    MB_D_FF_Float_147_183_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR147_183Output, Multiplier147WeightOutput);

    InputIEEE_Float_147_183: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier147WeightOutput, flopocoMultiplier147WeightOutput);

    MB_D_FF_Float_147_183_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier147WeightOutput, flopocoMultiplier147WeightInput);

    MB_D_FF_Float_Adder12_Input1_36_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier147_Output_183, mb_D_FFAdder12_Input1_36_0Output);

    MB_D_FF_Float_36_184_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder12_Input1_36_0Output, mb_D_FF36_184AugendStage1Output);

    MB_D_FF_Float_36_184_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF36_184AugendStage1Output, mb_D_FF36_184AugendStage2Output);

    Adder_Float_36: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF36_184AugendStage2Output, mb_D_FF36_184AddendStage2Output, Adder36_Output_184);

    MB_D_FF_Float_Adder12_Input2_36_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier142_Output_177, mb_D_FFAdder12_Input2_36_0Output);

    MB_D_FF_Float_36_184_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder12_Input2_36_0Output, mb_D_FF36_184AddendStage1Output);

    MB_D_FF_Float_36_184_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF36_184AddendStage1Output, mb_D_FF36_184AddendStage2Output);

    MB_D_FF_Float_Multiplier11_Input1_148_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder36_Output_184, mb_D_FFMultiplier11_Input1_148_0Output);

    MB_D_FF_Float_148_185_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier11_Input1_148_0Output, mb_D_FF148_185MultiplicandStage1Output);

    MB_D_FF_Float_148_185_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF148_185MultiplicandStage1Output, mb_D_FF148_185MultiplicandStage2Output);

    Multiplier_Float_148: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF148_185MultiplicandStage2Output, mb_D_FF148_185MultiplierStage2Output, Multiplier148_Output_185);

    MB_D_FF_Float_Multiplier11_Input2_148_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier137_Output_171, mb_D_FFMultiplier11_Input2_148_0Output);

    MB_D_FF_Float_148_185_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier11_Input2_148_0Output, mb_D_FF148_185MultiplierStage1Output);

    MB_D_FF_Float_148_185_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF148_185MultiplierStage1Output, mb_D_FF148_185MultiplierStage2Output);

    MB_D_FF_Float_Multiplier14_164_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier119_Output_147, mb_D_FFMultiplier14_164_0Output);

    MB_D_FF_Float_164_206_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier14_164_0Output, mb_D_FF164_206MultiplierStage1Output);

    MB_D_FF_Float_164_206_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF164_206MultiplierStage1Output, mb_D_FF164_206MultiplierStage2Output);

    Multiplier_Float_164: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF164_206MultiplierStage2Output, flopocoMultiplier164WeightInput, Multiplier164_Output_206);

    MBRightSHR_Float_164_206: entity work.MBRightSHR(rtl)
    GENERIC MAP (89, NumberOfBits)
    PORT MAP (clk, rst, Multiplier164Weight, mbRightSHR164_206Output);

    MB_D_FF_Float_164_206_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR164_206Output, Multiplier164WeightOutput);

    InputIEEE_Float_164_206: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier164WeightOutput, flopocoMultiplier164WeightOutput);

    MB_D_FF_Float_164_206_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier164WeightOutput, flopocoMultiplier164WeightInput);

    MB_D_FF_Float_Multiplier14_180_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier135_Output_168, mb_D_FFMultiplier14_180_0Output);

    MB_D_FF_Float_180_227_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier14_180_0Output, mb_D_FF180_227MultiplierStage1Output);

    MB_D_FF_Float_180_227_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF180_227MultiplierStage1Output, mb_D_FF180_227MultiplierStage2Output);

    Multiplier_Float_180: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF180_227MultiplierStage2Output, flopocoMultiplier180WeightInput, Multiplier180_Output_227);

    MBRightSHR_Float_180_227: entity work.MBRightSHR(rtl)
    GENERIC MAP (89, NumberOfBits)
    PORT MAP (clk, rst, Multiplier180Weight, mbRightSHR180_227Output);

    MB_D_FF_Float_180_227_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR180_227Output, Multiplier180WeightOutput);

    InputIEEE_Float_180_227: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier180WeightOutput, flopocoMultiplier180WeightOutput);

    MB_D_FF_Float_180_227_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier180WeightOutput, flopocoMultiplier180WeightInput);

    MB_D_FF_Float_Adder13_Input1_47_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier180_Output_227, mb_D_FFAdder13_Input1_47_0Output);

    MB_D_FF_Float_47_228_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder13_Input1_47_0Output, mb_D_FF47_228AugendStage1Output);

    MB_D_FF_Float_47_228_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF47_228AugendStage1Output, mb_D_FF47_228AugendStage2Output);

    Adder_Float_47: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF47_228AugendStage2Output, mb_D_FF47_228AddendStage2Output, Adder47_Output_228);

    MB_D_FF_Float_Adder13_Input2_47_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier164_Output_206, mb_D_FFAdder13_Input2_47_0Output);

    MB_D_FF_Float_47_228_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder13_Input2_47_0Output, mb_D_FF47_228AddendStage1Output);

    MB_D_FF_Float_47_228_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF47_228AddendStage1Output, mb_D_FF47_228AddendStage2Output);

    MB_D_FF_Float_Multiplier12_181_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder47_Output_228, mb_D_FFMultiplier12_181_0Output);

    MB_D_FF_Float_181_229_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier12_181_0Output, mb_D_FF181_229MultiplierStage1Output);

    MB_D_FF_Float_181_229_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF181_229MultiplierStage1Output, mb_D_FF181_229MultiplierStage2Output);

    Multiplier_Float_181: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF181_229MultiplierStage2Output, mb_D_FF181_229MultiplicandStage2Output, Multiplier181_Output_229);

    MBRightSHR_Float_181_229: entity work.MBRightSHR(rtl)
    GENERIC MAP (121, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR181_229Input, mbRightSHR181_229Output);

    MB_D_FF_Float_181_229_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR181_229Output, mb_D_FF181_229MultiplicandStage1Output);

    MB_D_FF_Float_181_229_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF181_229MultiplicandStage1Output, mb_D_FF181_229MultiplicandStage2Output);

    MBRightSHR_Float_182_Input1230: entity work.MBRightSHR(rtl)
    GENERIC MAP (50, NumberOfBits)
    PORT MAP (clk, rst, Multiplier182Weight, mbRightSHR182_Input1_230Output);

    MB_D_FF_Float_182_230_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR182_Input1_230Output, Multiplier182WeightOutput);

    InputIEEE_Float_182_230: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier182WeightOutput, flopocoMultiplier182WeightOutput);

    MB_D_FF_Float_182_230_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier182WeightOutput, flopocoMultiplier182WeightInput);

    Multiplier_Float_182: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier182WeightInput, mb_D_FF182_230MultiplierStage2Output, Multiplier182_Output_230);

    MBRightSHR_Float_182_Input2_230: entity work.MBRightSHR(rtl)
    GENERIC MAP (50, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR182_Input2_230Input, mbRightSHR182_Input2_230Output);

    MB_D_FF_Float_182_230_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR182_Input2_230Output, mb_D_FF182_230MultiplierStage1Output);

    MB_D_FF_Float_182_230_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF182_230MultiplierStage1Output, mb_D_FF182_230MultiplierStage2Output);

    MBRightSHR_Float_183_Input1231: entity work.MBRightSHR(rtl)
    GENERIC MAP (50, NumberOfBits)
    PORT MAP (clk, rst, Multiplier183Weight, mbRightSHR183_Input1_231Output);

    MB_D_FF_Float_183_231_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR183_Input1_231Output, Multiplier183WeightOutput);

    InputIEEE_Float_183_231: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier183WeightOutput, flopocoMultiplier183WeightOutput);

    MB_D_FF_Float_183_231_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier183WeightOutput, flopocoMultiplier183WeightInput);

    Multiplier_Float_183: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier183WeightInput, mb_D_FF183_231MultiplierStage2Output, Multiplier183_Output_231);

    MBRightSHR_Float_183_Input2_231: entity work.MBRightSHR(rtl)
    GENERIC MAP (50, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR183_Input2_231Input, mbRightSHR183_Input2_231Output);

    MB_D_FF_Float_183_231_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR183_Input2_231Output, mb_D_FF183_231MultiplierStage1Output);

    MB_D_FF_Float_183_231_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF183_231MultiplierStage1Output, mb_D_FF183_231MultiplierStage2Output);

    MB_D_FF_Float_Adder16_Input1_48_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier183_Output_231, mb_D_FFAdder16_Input1_48_0Output);

    MB_D_FF_Float_48_232_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder16_Input1_48_0Output, mb_D_FF48_232AugendStage1Output);

    MB_D_FF_Float_48_232_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF48_232AugendStage1Output, mb_D_FF48_232AugendStage2Output);

    Adder_Float_48: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF48_232AugendStage2Output, mb_D_FF48_232AddendStage2Output, Adder48_Output_232);

    MB_D_FF_Float_Adder16_Input2_48_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier182_Output_230, mb_D_FFAdder16_Input2_48_0Output);

    MB_D_FF_Float_48_232_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder16_Input2_48_0Output, mb_D_FF48_232AddendStage1Output);

    MB_D_FF_Float_48_232_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF48_232AddendStage1Output, mb_D_FF48_232AddendStage2Output);

    MB_D_FF_Float_Multiplier15_184_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder48_Output_232, mb_D_FFMultiplier15_184_0Output);

    MB_D_FF_Float_184_233_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier15_184_0Output, mb_D_FF184_233MultiplierStage1Output);

    MB_D_FF_Float_184_233_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF184_233MultiplierStage1Output, mb_D_FF184_233MultiplierStage2Output);

    Multiplier_Float_184: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF184_233MultiplierStage2Output, mb_D_FF184_233MultiplicandStage2Output, Multiplier184_Output_233);

    MBRightSHR_Float_184_233: entity work.MBRightSHR(rtl)
    GENERIC MAP (82, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR184_233Input, mbRightSHR184_233Output);

    MB_D_FF_Float_184_233_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR184_233Output, mb_D_FF184_233MultiplicandStage1Output);

    MB_D_FF_Float_184_233_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF184_233MultiplicandStage1Output, mb_D_FF184_233MultiplicandStage2Output);

    MB_D_FF_Float_Multiplier14_185_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier184_Output_233, mb_D_FFMultiplier14_185_0Output);

    MB_D_FF_Float_185_234_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier14_185_0Output, mb_D_FF185_234MultiplierStage1Output);

    MB_D_FF_Float_185_234_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF185_234MultiplierStage1Output, mb_D_FF185_234MultiplierStage2Output);

    Multiplier_Float_185: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF185_234MultiplierStage2Output, flopocoMultiplier185WeightInput, Multiplier185_Output_234);

    MBRightSHR_Float_185_234: entity work.MBRightSHR(rtl)
    GENERIC MAP (89, NumberOfBits)
    PORT MAP (clk, rst, Multiplier185Weight, mbRightSHR185_234Output);

    MB_D_FF_Float_185_234_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR185_234Output, Multiplier185WeightOutput);

    InputIEEE_Float_185_234: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier185WeightOutput, flopocoMultiplier185WeightOutput);

    MB_D_FF_Float_185_234_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier185WeightOutput, flopocoMultiplier185WeightInput);

    MB_D_FF_Float_Multiplier13_186_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier185_Output_234, mb_D_FFMultiplier13_186_0Output);

    MB_D_FF_Float_186_235_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier13_186_0Output, mb_D_FF186_235MultiplierStage1Output);

    MB_D_FF_Float_186_235_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF186_235MultiplierStage1Output, mb_D_FF186_235MultiplierStage2Output);

    Multiplier_Float_186: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF186_235MultiplierStage2Output, flopocoMultiplier186WeightInput, Multiplier186_Output_235);

    MBRightSHR_Float_186_235: entity work.MBRightSHR(rtl)
    GENERIC MAP (96, NumberOfBits)
    PORT MAP (clk, rst, Multiplier186Weight, mbRightSHR186_235Output);

    MB_D_FF_Float_186_235_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR186_235Output, Multiplier186WeightOutput);

    InputIEEE_Float_186_235: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier186WeightOutput, flopocoMultiplier186WeightOutput);

    MB_D_FF_Float_186_235_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier186WeightOutput, flopocoMultiplier186WeightInput);

    MBRightSHR_Float_187_Input1236: entity work.MBRightSHR(rtl)
    GENERIC MAP (50, NumberOfBits)
    PORT MAP (clk, rst, Multiplier187Weight, mbRightSHR187_Input1_236Output);

    MB_D_FF_Float_187_236_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR187_Input1_236Output, Multiplier187WeightOutput);

    InputIEEE_Float_187_236: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier187WeightOutput, flopocoMultiplier187WeightOutput);

    MB_D_FF_Float_187_236_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier187WeightOutput, flopocoMultiplier187WeightInput);

    Multiplier_Float_187: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier187WeightInput, mb_D_FF187_236MultiplierStage2Output, Multiplier187_Output_236);

    MBRightSHR_Float_187_Input2_236: entity work.MBRightSHR(rtl)
    GENERIC MAP (50, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR187_Input2_236Input, mbRightSHR187_Input2_236Output);

    MB_D_FF_Float_187_236_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR187_Input2_236Output, mb_D_FF187_236MultiplierStage1Output);

    MB_D_FF_Float_187_236_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF187_236MultiplierStage1Output, mb_D_FF187_236MultiplierStage2Output);

    MBRightSHR_Float_188_Input1237: entity work.MBRightSHR(rtl)
    GENERIC MAP (50, NumberOfBits)
    PORT MAP (clk, rst, Multiplier188Weight, mbRightSHR188_Input1_237Output);

    MB_D_FF_Float_188_237_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR188_Input1_237Output, Multiplier188WeightOutput);

    InputIEEE_Float_188_237: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier188WeightOutput, flopocoMultiplier188WeightOutput);

    MB_D_FF_Float_188_237_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier188WeightOutput, flopocoMultiplier188WeightInput);

    Multiplier_Float_188: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier188WeightInput, mb_D_FF188_237MultiplierStage2Output, Multiplier188_Output_237);

    MBRightSHR_Float_188_Input2_237: entity work.MBRightSHR(rtl)
    GENERIC MAP (50, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR188_Input2_237Input, mbRightSHR188_Input2_237Output);

    MB_D_FF_Float_188_237_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR188_Input2_237Output, mb_D_FF188_237MultiplierStage1Output);

    MB_D_FF_Float_188_237_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF188_237MultiplierStage1Output, mb_D_FF188_237MultiplierStage2Output);

    MB_D_FF_Float_Adder16_Input1_49_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier188_Output_237, mb_D_FFAdder16_Input1_49_0Output);

    MB_D_FF_Float_49_238_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder16_Input1_49_0Output, mb_D_FF49_238AugendStage1Output);

    MB_D_FF_Float_49_238_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF49_238AugendStage1Output, mb_D_FF49_238AugendStage2Output);

    Adder_Float_49: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF49_238AugendStage2Output, mb_D_FF49_238AddendStage2Output, Adder49_Output_238);

    MB_D_FF_Float_Adder16_Input2_49_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier187_Output_236, mb_D_FFAdder16_Input2_49_0Output);

    MB_D_FF_Float_49_238_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder16_Input2_49_0Output, mb_D_FF49_238AddendStage1Output);

    MB_D_FF_Float_49_238_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF49_238AddendStage1Output, mb_D_FF49_238AddendStage2Output);

    MB_D_FF_Float_Multiplier15_189_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder49_Output_238, mb_D_FFMultiplier15_189_0Output);

    MB_D_FF_Float_189_239_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier15_189_0Output, mb_D_FF189_239MultiplierStage1Output);

    MB_D_FF_Float_189_239_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF189_239MultiplierStage1Output, mb_D_FF189_239MultiplierStage2Output);

    Multiplier_Float_189: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF189_239MultiplierStage2Output, mb_D_FF189_239MultiplicandStage2Output, Multiplier189_Output_239);

    MBRightSHR_Float_189_239: entity work.MBRightSHR(rtl)
    GENERIC MAP (82, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR189_239Input, mbRightSHR189_239Output);

    MB_D_FF_Float_189_239_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR189_239Output, mb_D_FF189_239MultiplicandStage1Output);

    MB_D_FF_Float_189_239_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF189_239MultiplicandStage1Output, mb_D_FF189_239MultiplicandStage2Output);

    MB_D_FF_Float_Multiplier14_190_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier189_Output_239, mb_D_FFMultiplier14_190_0Output);

    MB_D_FF_Float_190_240_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier14_190_0Output, mb_D_FF190_240MultiplierStage1Output);

    MB_D_FF_Float_190_240_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF190_240MultiplierStage1Output, mb_D_FF190_240MultiplierStage2Output);

    Multiplier_Float_190: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF190_240MultiplierStage2Output, flopocoMultiplier190WeightInput, Multiplier190_Output_240);

    MBRightSHR_Float_190_240: entity work.MBRightSHR(rtl)
    GENERIC MAP (89, NumberOfBits)
    PORT MAP (clk, rst, Multiplier190Weight, mbRightSHR190_240Output);

    MB_D_FF_Float_190_240_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR190_240Output, Multiplier190WeightOutput);

    InputIEEE_Float_190_240: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier190WeightOutput, flopocoMultiplier190WeightOutput);

    MB_D_FF_Float_190_240_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier190WeightOutput, flopocoMultiplier190WeightInput);

    MB_D_FF_Float_Multiplier13_191_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier190_Output_240, mb_D_FFMultiplier13_191_0Output);

    MB_D_FF_Float_191_241_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier13_191_0Output, mb_D_FF191_241MultiplierStage1Output);

    MB_D_FF_Float_191_241_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF191_241MultiplierStage1Output, mb_D_FF191_241MultiplierStage2Output);

    Multiplier_Float_191: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF191_241MultiplierStage2Output, flopocoMultiplier191WeightInput, Multiplier191_Output_241);

    MBRightSHR_Float_191_241: entity work.MBRightSHR(rtl)
    GENERIC MAP (96, NumberOfBits)
    PORT MAP (clk, rst, Multiplier191Weight, mbRightSHR191_241Output);

    MB_D_FF_Float_191_241_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR191_241Output, Multiplier191WeightOutput);

    InputIEEE_Float_191_241: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier191WeightOutput, flopocoMultiplier191WeightOutput);

    MB_D_FF_Float_191_241_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier191WeightOutput, flopocoMultiplier191WeightInput);

    MB_D_FF_Float_Adder12_Input1_50_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier191_Output_241, mb_D_FFAdder12_Input1_50_0Output);

    MB_D_FF_Float_50_242_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder12_Input1_50_0Output, mb_D_FF50_242AugendStage1Output);

    MB_D_FF_Float_50_242_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF50_242AugendStage1Output, mb_D_FF50_242AugendStage2Output);

    Adder_Float_50: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF50_242AugendStage2Output, mb_D_FF50_242AddendStage2Output, Adder50_Output_242);

    MB_D_FF_Float_Adder12_Input2_50_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier186_Output_235, mb_D_FFAdder12_Input2_50_0Output);

    MB_D_FF_Float_50_242_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder12_Input2_50_0Output, mb_D_FF50_242AddendStage1Output);

    MB_D_FF_Float_50_242_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF50_242AddendStage1Output, mb_D_FF50_242AddendStage2Output);

    MB_D_FF_Float_Multiplier11_Input1_192_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder50_Output_242, mb_D_FFMultiplier11_Input1_192_0Output);

    MB_D_FF_Float_192_243_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier11_Input1_192_0Output, mb_D_FF192_243MultiplicandStage1Output);

    MB_D_FF_Float_192_243_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF192_243MultiplicandStage1Output, mb_D_FF192_243MultiplicandStage2Output);

    Multiplier_Float_192: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF192_243MultiplicandStage2Output, mb_D_FF192_243MultiplierStage2Output, Multiplier192_Output_243);

    MB_D_FF_Float_Multiplier11_Input2_192_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier181_Output_229, mb_D_FFMultiplier11_Input2_192_0Output);

    MB_D_FF_Float_192_243_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier11_Input2_192_0Output, mb_D_FF192_243MultiplierStage1Output);

    MB_D_FF_Float_192_243_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF192_243MultiplierStage1Output, mb_D_FF192_243MultiplierStage2Output);

    MB_D_FF_Float_Adder10_Input1_51_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier192_Output_243, mb_D_FFAdder10_Input1_51_0Output);

    MB_D_FF_Float_51_244_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder10_Input1_51_0Output, mb_D_FF51_244AugendStage1Output);

    MB_D_FF_Float_51_244_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF51_244AugendStage1Output, mb_D_FF51_244AugendStage2Output);

    Adder_Float_51: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF51_244AugendStage2Output, mb_D_FF51_244AddendStage2Output, Adder51_Output_244);

    MB_D_FF_Float_Adder10_Input2_51_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier148_Output_185, mb_D_FFAdder10_Input2_51_0Output);

    MB_D_FF_Float_51_244_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder10_Input2_51_0Output, mb_D_FF51_244AddendStage1Output);

    MB_D_FF_Float_51_244_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF51_244AddendStage1Output, mb_D_FF51_244AddendStage2Output);

    MB_D_FF_Float_Multiplier9_193_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder51_Output_244, mb_D_FFMultiplier9_193_0Output);

    MB_D_FF_Float_193_245_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier9_193_0Output, mb_D_FF193_245MultiplierStage1Output);

    MB_D_FF_Float_193_245_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF193_245MultiplierStage1Output, mb_D_FF193_245MultiplierStage2Output);

    Multiplier_Float_193: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF193_245MultiplierStage2Output, mb_D_FF193_245MultiplicandStage2Output, Multiplier193_Output_245);

    MBRightSHR_Float_193_245: entity work.MBRightSHR(rtl)
    GENERIC MAP (160, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR193_245Input, mbRightSHR193_245Output);

    MB_D_FF_Float_193_245_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR193_245Output, mb_D_FF193_245MultiplicandStage1Output);

    MB_D_FF_Float_193_245_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF193_245MultiplicandStage1Output, mb_D_FF193_245MultiplicandStage2Output);

    MB_D_FF_Float_Multiplier8_194_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier193_Output_245, mb_D_FFMultiplier8_194_0Output);

    MB_D_FF_Float_194_246_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier8_194_0Output, mb_D_FF194_246MultiplierStage1Output);

    MB_D_FF_Float_194_246_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF194_246MultiplierStage1Output, mb_D_FF194_246MultiplierStage2Output);

    Multiplier_Float_194: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF194_246MultiplierStage2Output, flopocoMultiplier194WeightInput, Multiplier194_Output_246);

    MBRightSHR_Float_194_246: entity work.MBRightSHR(rtl)
    GENERIC MAP (167, NumberOfBits)
    PORT MAP (clk, rst, Multiplier194Weight, mbRightSHR194_246Output);

    MB_D_FF_Float_194_246_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR194_246Output, Multiplier194WeightOutput);

    InputIEEE_Float_194_246: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier194WeightOutput, flopocoMultiplier194WeightOutput);

    MB_D_FF_Float_194_246_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier194WeightOutput, flopocoMultiplier194WeightInput);

    MBRightSHR_Float_199_Input1252: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits)
    PORT MAP (clk, rst, Multiplier199Weight, mbRightSHR199_Input1_252Output);

    MB_D_FF_Float_199_252_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR199_Input1_252Output, Multiplier199WeightOutput);

    InputIEEE_Float_199_252: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier199WeightOutput, flopocoMultiplier199WeightOutput);

    MB_D_FF_Float_199_252_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier199WeightOutput, flopocoMultiplier199WeightInput);

    Multiplier_Float_199: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier199WeightInput, mb_D_FF199_252MultiplierStage2Output, Multiplier199_Output_252);

    MBRightSHR_Float_199_Input2_252: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR199_Input2_252Input, mbRightSHR199_Input2_252Output);

    MB_D_FF_Float_199_252_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR199_Input2_252Output, mb_D_FF199_252MultiplierStage1Output);

    MB_D_FF_Float_199_252_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF199_252MultiplierStage1Output, mb_D_FF199_252MultiplierStage2Output);

    MBRightSHR_Float_200_Input1253: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits)
    PORT MAP (clk, rst, Multiplier200Weight, mbRightSHR200_Input1_253Output);

    MB_D_FF_Float_200_253_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR200_Input1_253Output, Multiplier200WeightOutput);

    InputIEEE_Float_200_253: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier200WeightOutput, flopocoMultiplier200WeightOutput);

    MB_D_FF_Float_200_253_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier200WeightOutput, flopocoMultiplier200WeightInput);

    Multiplier_Float_200: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier200WeightInput, mb_D_FF200_253MultiplierStage2Output, Multiplier200_Output_253);

    MBRightSHR_Float_200_Input2_253: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR200_Input2_253Input, mbRightSHR200_Input2_253Output);

    MB_D_FF_Float_200_253_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR200_Input2_253Output, mb_D_FF200_253MultiplierStage1Output);

    MB_D_FF_Float_200_253_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF200_253MultiplierStage1Output, mb_D_FF200_253MultiplierStage2Output);

    MB_D_FF_Float_Adder18_Input1_53_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier200_Output_253, mb_D_FFAdder18_Input1_53_0Output);

    MB_D_FF_Float_53_254_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder18_Input1_53_0Output, mb_D_FF53_254AugendStage1Output);

    MB_D_FF_Float_53_254_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF53_254AugendStage1Output, mb_D_FF53_254AugendStage2Output);

    Adder_Float_53: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF53_254AugendStage2Output, mb_D_FF53_254AddendStage2Output, Adder53_Output_254);

    MB_D_FF_Float_Adder18_Input2_53_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier199_Output_252, mb_D_FFAdder18_Input2_53_0Output);

    MB_D_FF_Float_53_254_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder18_Input2_53_0Output, mb_D_FF53_254AddendStage1Output);

    MB_D_FF_Float_53_254_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF53_254AddendStage1Output, mb_D_FF53_254AddendStage2Output);

    MB_D_FF_Float_Multiplier17_Input1_201_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder53_Output_254, mb_D_FFMultiplier17_Input1_201_0Output);

    MB_D_FF_Float_201_255_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier17_Input1_201_0Output, mb_D_FF201_255MultiplicandStage1Output);

    MB_D_FF_Float_201_255_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF201_255MultiplicandStage1Output, mb_D_FF201_255MultiplicandStage2Output);

    Multiplier_Float_201: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF201_255MultiplicandStage2Output, mb_D_FF201_255MultiplierStage2Output, Multiplier201_Output_255);

    MB_D_FF_Float_Multiplier17_Input2_201_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier108_Output_132, mb_D_FFMultiplier17_Input2_201_0Output);

    MB_D_FF_Float_201_255_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier17_Input2_201_0Output, mb_D_FF201_255MultiplierStage1Output);

    MB_D_FF_Float_201_255_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF201_255MultiplierStage1Output, mb_D_FF201_255MultiplierStage2Output);

    MBRightSHR_Float_206_Input1261: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits)
    PORT MAP (clk, rst, Multiplier206Weight, mbRightSHR206_Input1_261Output);

    MB_D_FF_Float_206_261_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR206_Input1_261Output, Multiplier206WeightOutput);

    InputIEEE_Float_206_261: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier206WeightOutput, flopocoMultiplier206WeightOutput);

    MB_D_FF_Float_206_261_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier206WeightOutput, flopocoMultiplier206WeightInput);

    Multiplier_Float_206: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier206WeightInput, mb_D_FF206_261MultiplierStage2Output, Multiplier206_Output_261);

    MBRightSHR_Float_206_Input2_261: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR206_Input2_261Input, mbRightSHR206_Input2_261Output);

    MB_D_FF_Float_206_261_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR206_Input2_261Output, mb_D_FF206_261MultiplierStage1Output);

    MB_D_FF_Float_206_261_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF206_261MultiplierStage1Output, mb_D_FF206_261MultiplierStage2Output);

    MBRightSHR_Float_207_Input1262: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits)
    PORT MAP (clk, rst, Multiplier207Weight, mbRightSHR207_Input1_262Output);

    MB_D_FF_Float_207_262_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR207_Input1_262Output, Multiplier207WeightOutput);

    InputIEEE_Float_207_262: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier207WeightOutput, flopocoMultiplier207WeightOutput);

    MB_D_FF_Float_207_262_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier207WeightOutput, flopocoMultiplier207WeightInput);

    Multiplier_Float_207: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier207WeightInput, mb_D_FF207_262MultiplierStage2Output, Multiplier207_Output_262);

    MBRightSHR_Float_207_Input2_262: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR207_Input2_262Input, mbRightSHR207_Input2_262Output);

    MB_D_FF_Float_207_262_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR207_Input2_262Output, mb_D_FF207_262MultiplierStage1Output);

    MB_D_FF_Float_207_262_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF207_262MultiplierStage1Output, mb_D_FF207_262MultiplierStage2Output);

    MB_D_FF_Float_Adder18_Input1_55_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier207_Output_262, mb_D_FFAdder18_Input1_55_0Output);

    MB_D_FF_Float_55_263_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder18_Input1_55_0Output, mb_D_FF55_263AugendStage1Output);

    MB_D_FF_Float_55_263_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF55_263AugendStage1Output, mb_D_FF55_263AugendStage2Output);

    Adder_Float_55: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF55_263AugendStage2Output, mb_D_FF55_263AddendStage2Output, Adder55_Output_263);

    MB_D_FF_Float_Adder18_Input2_55_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier206_Output_261, mb_D_FFAdder18_Input2_55_0Output);

    MB_D_FF_Float_55_263_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder18_Input2_55_0Output, mb_D_FF55_263AddendStage1Output);

    MB_D_FF_Float_55_263_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF55_263AddendStage1Output, mb_D_FF55_263AddendStage2Output);

    MB_D_FF_Float_Multiplier17_Input1_208_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder55_Output_263, mb_D_FFMultiplier17_Input1_208_0Output);

    MB_D_FF_Float_208_264_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier17_Input1_208_0Output, mb_D_FF208_264MultiplicandStage1Output);

    MB_D_FF_Float_208_264_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF208_264MultiplicandStage1Output, mb_D_FF208_264MultiplicandStage2Output);

    Multiplier_Float_208: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF208_264MultiplicandStage2Output, mb_D_FF208_264MultiplierStage2Output, Multiplier208_Output_264);

    MB_D_FF_Float_Multiplier17_Input2_208_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier115_Output_141, mb_D_FFMultiplier17_Input2_208_0Output);

    MB_D_FF_Float_208_264_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier17_Input2_208_0Output, mb_D_FF208_264MultiplierStage1Output);

    MB_D_FF_Float_208_264_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF208_264MultiplierStage1Output, mb_D_FF208_264MultiplierStage2Output);

    MB_D_FF_Float_Adder16_Input1_56_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier208_Output_264, mb_D_FFAdder16_Input1_56_0Output);

    MB_D_FF_Float_56_265_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder16_Input1_56_0Output, mb_D_FF56_265AugendStage1Output);

    MB_D_FF_Float_56_265_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF56_265AugendStage1Output, mb_D_FF56_265AugendStage2Output);

    Adder_Float_56: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF56_265AugendStage2Output, mb_D_FF56_265AddendStage2Output, Adder56_Output_265);

    MB_D_FF_Float_Adder16_Input2_56_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier201_Output_255, mb_D_FFAdder16_Input2_56_0Output);

    MB_D_FF_Float_56_265_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder16_Input2_56_0Output, mb_D_FF56_265AddendStage1Output);

    MB_D_FF_Float_56_265_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF56_265AddendStage1Output, mb_D_FF56_265AddendStage2Output);

    MB_D_FF_Float_Multiplier15_209_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder56_Output_265, mb_D_FFMultiplier15_209_0Output);

    MB_D_FF_Float_209_266_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier15_209_0Output, mb_D_FF209_266MultiplierStage1Output);

    MB_D_FF_Float_209_266_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF209_266MultiplierStage1Output, mb_D_FF209_266MultiplierStage2Output);

    Multiplier_Float_209: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF209_266MultiplierStage2Output, mb_D_FF209_266MultiplicandStage2Output, Multiplier209_Output_266);

    MBRightSHR_Float_209_266: entity work.MBRightSHR(rtl)
    GENERIC MAP (82, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR209_266Input, mbRightSHR209_266Output);

    MB_D_FF_Float_209_266_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR209_266Output, mb_D_FF209_266MultiplicandStage1Output);

    MB_D_FF_Float_209_266_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF209_266MultiplicandStage1Output, mb_D_FF209_266MultiplicandStage2Output);

    MB_D_FF_Float_Multiplier14_210_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier209_Output_266, mb_D_FFMultiplier14_210_0Output);

    MB_D_FF_Float_210_267_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier14_210_0Output, mb_D_FF210_267MultiplierStage1Output);

    MB_D_FF_Float_210_267_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF210_267MultiplierStage1Output, mb_D_FF210_267MultiplierStage2Output);

    Multiplier_Float_210: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF210_267MultiplierStage2Output, flopocoMultiplier210WeightInput, Multiplier210_Output_267);

    MBRightSHR_Float_210_267: entity work.MBRightSHR(rtl)
    GENERIC MAP (89, NumberOfBits)
    PORT MAP (clk, rst, Multiplier210Weight, mbRightSHR210_267Output);

    MB_D_FF_Float_210_267_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR210_267Output, Multiplier210WeightOutput);

    InputIEEE_Float_210_267: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier210WeightOutput, flopocoMultiplier210WeightOutput);

    MB_D_FF_Float_210_267_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier210WeightOutput, flopocoMultiplier210WeightInput);

    MBRightSHR_Float_215_Input1273: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits)
    PORT MAP (clk, rst, Multiplier215Weight, mbRightSHR215_Input1_273Output);

    MB_D_FF_Float_215_273_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR215_Input1_273Output, Multiplier215WeightOutput);

    InputIEEE_Float_215_273: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier215WeightOutput, flopocoMultiplier215WeightOutput);

    MB_D_FF_Float_215_273_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier215WeightOutput, flopocoMultiplier215WeightInput);

    Multiplier_Float_215: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier215WeightInput, mb_D_FF215_273MultiplierStage2Output, Multiplier215_Output_273);

    MBRightSHR_Float_215_Input2_273: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR215_Input2_273Input, mbRightSHR215_Input2_273Output);

    MB_D_FF_Float_215_273_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR215_Input2_273Output, mb_D_FF215_273MultiplierStage1Output);

    MB_D_FF_Float_215_273_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF215_273MultiplierStage1Output, mb_D_FF215_273MultiplierStage2Output);

    MBRightSHR_Float_216_Input1274: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits)
    PORT MAP (clk, rst, Multiplier216Weight, mbRightSHR216_Input1_274Output);

    MB_D_FF_Float_216_274_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR216_Input1_274Output, Multiplier216WeightOutput);

    InputIEEE_Float_216_274: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier216WeightOutput, flopocoMultiplier216WeightOutput);

    MB_D_FF_Float_216_274_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier216WeightOutput, flopocoMultiplier216WeightInput);

    Multiplier_Float_216: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier216WeightInput, mb_D_FF216_274MultiplierStage2Output, Multiplier216_Output_274);

    MBRightSHR_Float_216_Input2_274: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR216_Input2_274Input, mbRightSHR216_Input2_274Output);

    MB_D_FF_Float_216_274_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR216_Input2_274Output, mb_D_FF216_274MultiplierStage1Output);

    MB_D_FF_Float_216_274_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF216_274MultiplierStage1Output, mb_D_FF216_274MultiplierStage2Output);

    MB_D_FF_Float_Adder18_Input1_58_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier216_Output_274, mb_D_FFAdder18_Input1_58_0Output);

    MB_D_FF_Float_58_275_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder18_Input1_58_0Output, mb_D_FF58_275AugendStage1Output);

    MB_D_FF_Float_58_275_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF58_275AugendStage1Output, mb_D_FF58_275AugendStage2Output);

    Adder_Float_58: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF58_275AugendStage2Output, mb_D_FF58_275AddendStage2Output, Adder58_Output_275);

    MB_D_FF_Float_Adder18_Input2_58_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier215_Output_273, mb_D_FFAdder18_Input2_58_0Output);

    MB_D_FF_Float_58_275_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder18_Input2_58_0Output, mb_D_FF58_275AddendStage1Output);

    MB_D_FF_Float_58_275_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF58_275AddendStage1Output, mb_D_FF58_275AddendStage2Output);

    MB_D_FF_Float_Multiplier17_Input1_217_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder58_Output_275, mb_D_FFMultiplier17_Input1_217_0Output);

    MB_D_FF_Float_217_276_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier17_Input1_217_0Output, mb_D_FF217_276MultiplicandStage1Output);

    MB_D_FF_Float_217_276_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF217_276MultiplicandStage1Output, mb_D_FF217_276MultiplicandStage2Output);

    Multiplier_Float_217: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF217_276MultiplicandStage2Output, mb_D_FF217_276MultiplierStage2Output, Multiplier217_Output_276);

    MB_D_FF_Float_Multiplier17_Input2_217_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier124_Output_153, mb_D_FFMultiplier17_Input2_217_0Output);

    MB_D_FF_Float_217_276_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier17_Input2_217_0Output, mb_D_FF217_276MultiplierStage1Output);

    MB_D_FF_Float_217_276_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF217_276MultiplierStage1Output, mb_D_FF217_276MultiplierStage2Output);

    MBRightSHR_Float_222_Input1282: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits)
    PORT MAP (clk, rst, Multiplier222Weight, mbRightSHR222_Input1_282Output);

    MB_D_FF_Float_222_282_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR222_Input1_282Output, Multiplier222WeightOutput);

    InputIEEE_Float_222_282: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier222WeightOutput, flopocoMultiplier222WeightOutput);

    MB_D_FF_Float_222_282_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier222WeightOutput, flopocoMultiplier222WeightInput);

    Multiplier_Float_222: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier222WeightInput, mb_D_FF222_282MultiplierStage2Output, Multiplier222_Output_282);

    MBRightSHR_Float_222_Input2_282: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR222_Input2_282Input, mbRightSHR222_Input2_282Output);

    MB_D_FF_Float_222_282_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR222_Input2_282Output, mb_D_FF222_282MultiplierStage1Output);

    MB_D_FF_Float_222_282_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF222_282MultiplierStage1Output, mb_D_FF222_282MultiplierStage2Output);

    MBRightSHR_Float_223_Input1283: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits)
    PORT MAP (clk, rst, Multiplier223Weight, mbRightSHR223_Input1_283Output);

    MB_D_FF_Float_223_283_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR223_Input1_283Output, Multiplier223WeightOutput);

    InputIEEE_Float_223_283: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier223WeightOutput, flopocoMultiplier223WeightOutput);

    MB_D_FF_Float_223_283_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier223WeightOutput, flopocoMultiplier223WeightInput);

    Multiplier_Float_223: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier223WeightInput, mb_D_FF223_283MultiplierStage2Output, Multiplier223_Output_283);

    MBRightSHR_Float_223_Input2_283: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR223_Input2_283Input, mbRightSHR223_Input2_283Output);

    MB_D_FF_Float_223_283_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR223_Input2_283Output, mb_D_FF223_283MultiplierStage1Output);

    MB_D_FF_Float_223_283_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF223_283MultiplierStage1Output, mb_D_FF223_283MultiplierStage2Output);

    MB_D_FF_Float_Adder18_Input1_60_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier223_Output_283, mb_D_FFAdder18_Input1_60_0Output);

    MB_D_FF_Float_60_284_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder18_Input1_60_0Output, mb_D_FF60_284AugendStage1Output);

    MB_D_FF_Float_60_284_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF60_284AugendStage1Output, mb_D_FF60_284AugendStage2Output);

    Adder_Float_60: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF60_284AugendStage2Output, mb_D_FF60_284AddendStage2Output, Adder60_Output_284);

    MB_D_FF_Float_Adder18_Input2_60_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier222_Output_282, mb_D_FFAdder18_Input2_60_0Output);

    MB_D_FF_Float_60_284_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder18_Input2_60_0Output, mb_D_FF60_284AddendStage1Output);

    MB_D_FF_Float_60_284_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF60_284AddendStage1Output, mb_D_FF60_284AddendStage2Output);

    MB_D_FF_Float_Multiplier17_Input1_224_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder60_Output_284, mb_D_FFMultiplier17_Input1_224_0Output);

    MB_D_FF_Float_224_285_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier17_Input1_224_0Output, mb_D_FF224_285MultiplicandStage1Output);

    MB_D_FF_Float_224_285_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF224_285MultiplicandStage1Output, mb_D_FF224_285MultiplicandStage2Output);

    Multiplier_Float_224: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF224_285MultiplicandStage2Output, mb_D_FF224_285MultiplierStage2Output, Multiplier224_Output_285);

    MB_D_FF_Float_Multiplier17_Input2_224_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier131_Output_162, mb_D_FFMultiplier17_Input2_224_0Output);

    MB_D_FF_Float_224_285_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier17_Input2_224_0Output, mb_D_FF224_285MultiplierStage1Output);

    MB_D_FF_Float_224_285_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF224_285MultiplierStage1Output, mb_D_FF224_285MultiplierStage2Output);

    MB_D_FF_Float_Adder16_Input1_61_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier224_Output_285, mb_D_FFAdder16_Input1_61_0Output);

    MB_D_FF_Float_61_286_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder16_Input1_61_0Output, mb_D_FF61_286AugendStage1Output);

    MB_D_FF_Float_61_286_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF61_286AugendStage1Output, mb_D_FF61_286AugendStage2Output);

    Adder_Float_61: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF61_286AugendStage2Output, mb_D_FF61_286AddendStage2Output, Adder61_Output_286);

    MB_D_FF_Float_Adder16_Input2_61_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier217_Output_276, mb_D_FFAdder16_Input2_61_0Output);

    MB_D_FF_Float_61_286_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder16_Input2_61_0Output, mb_D_FF61_286AddendStage1Output);

    MB_D_FF_Float_61_286_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF61_286AddendStage1Output, mb_D_FF61_286AddendStage2Output);

    MB_D_FF_Float_Multiplier15_225_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder61_Output_286, mb_D_FFMultiplier15_225_0Output);

    MB_D_FF_Float_225_287_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier15_225_0Output, mb_D_FF225_287MultiplierStage1Output);

    MB_D_FF_Float_225_287_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF225_287MultiplierStage1Output, mb_D_FF225_287MultiplierStage2Output);

    Multiplier_Float_225: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF225_287MultiplierStage2Output, mb_D_FF225_287MultiplicandStage2Output, Multiplier225_Output_287);

    MBRightSHR_Float_225_287: entity work.MBRightSHR(rtl)
    GENERIC MAP (82, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR225_287Input, mbRightSHR225_287Output);

    MB_D_FF_Float_225_287_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR225_287Output, mb_D_FF225_287MultiplicandStage1Output);

    MB_D_FF_Float_225_287_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF225_287MultiplicandStage1Output, mb_D_FF225_287MultiplicandStage2Output);

    MB_D_FF_Float_Multiplier14_226_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier225_Output_287, mb_D_FFMultiplier14_226_0Output);

    MB_D_FF_Float_226_288_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier14_226_0Output, mb_D_FF226_288MultiplierStage1Output);

    MB_D_FF_Float_226_288_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF226_288MultiplierStage1Output, mb_D_FF226_288MultiplierStage2Output);

    Multiplier_Float_226: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF226_288MultiplierStage2Output, flopocoMultiplier226WeightInput, Multiplier226_Output_288);

    MBRightSHR_Float_226_288: entity work.MBRightSHR(rtl)
    GENERIC MAP (89, NumberOfBits)
    PORT MAP (clk, rst, Multiplier226Weight, mbRightSHR226_288Output);

    MB_D_FF_Float_226_288_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR226_288Output, Multiplier226WeightOutput);

    InputIEEE_Float_226_288: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier226WeightOutput, flopocoMultiplier226WeightOutput);

    MB_D_FF_Float_226_288_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier226WeightOutput, flopocoMultiplier226WeightInput);

    MB_D_FF_Float_Adder13_Input1_62_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier226_Output_288, mb_D_FFAdder13_Input1_62_0Output);

    MB_D_FF_Float_62_289_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder13_Input1_62_0Output, mb_D_FF62_289AugendStage1Output);

    MB_D_FF_Float_62_289_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF62_289AugendStage1Output, mb_D_FF62_289AugendStage2Output);

    Adder_Float_62: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF62_289AugendStage2Output, mb_D_FF62_289AddendStage2Output, Adder62_Output_289);

    MB_D_FF_Float_Adder13_Input2_62_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier210_Output_267, mb_D_FFAdder13_Input2_62_0Output);

    MB_D_FF_Float_62_289_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder13_Input2_62_0Output, mb_D_FF62_289AddendStage1Output);

    MB_D_FF_Float_62_289_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF62_289AddendStage1Output, mb_D_FF62_289AddendStage2Output);

    MB_D_FF_Float_Multiplier12_227_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder62_Output_289, mb_D_FFMultiplier12_227_0Output);

    MB_D_FF_Float_227_290_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier12_227_0Output, mb_D_FF227_290MultiplierStage1Output);

    MB_D_FF_Float_227_290_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF227_290MultiplierStage1Output, mb_D_FF227_290MultiplierStage2Output);

    Multiplier_Float_227: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF227_290MultiplierStage2Output, mb_D_FF227_290MultiplicandStage2Output, Multiplier227_Output_290);

    MBRightSHR_Float_227_290: entity work.MBRightSHR(rtl)
    GENERIC MAP (121, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR227_290Input, mbRightSHR227_290Output);

    MB_D_FF_Float_227_290_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR227_290Output, mb_D_FF227_290MultiplicandStage1Output);

    MB_D_FF_Float_227_290_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF227_290MultiplicandStage1Output, mb_D_FF227_290MultiplicandStage2Output);

    MB_D_FF_Float_Multiplier14_231_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier140_Output_175, mb_D_FFMultiplier14_231_0Output);

    MB_D_FF_Float_231_295_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier14_231_0Output, mb_D_FF231_295MultiplierStage1Output);

    MB_D_FF_Float_231_295_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF231_295MultiplierStage1Output, mb_D_FF231_295MultiplierStage2Output);

    Multiplier_Float_231: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF231_295MultiplierStage2Output, flopocoMultiplier231WeightInput, Multiplier231_Output_295);

    MBRightSHR_Float_231_295: entity work.MBRightSHR(rtl)
    GENERIC MAP (89, NumberOfBits)
    PORT MAP (clk, rst, Multiplier231Weight, mbRightSHR231_295Output);

    MB_D_FF_Float_231_295_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR231_295Output, Multiplier231WeightOutput);

    InputIEEE_Float_231_295: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier231WeightOutput, flopocoMultiplier231WeightOutput);

    MB_D_FF_Float_231_295_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier231WeightOutput, flopocoMultiplier231WeightInput);

    MB_D_FF_Float_Multiplier13_232_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier231_Output_295, mb_D_FFMultiplier13_232_0Output);

    MB_D_FF_Float_232_296_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier13_232_0Output, mb_D_FF232_296MultiplierStage1Output);

    MB_D_FF_Float_232_296_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF232_296MultiplierStage1Output, mb_D_FF232_296MultiplierStage2Output);

    Multiplier_Float_232: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF232_296MultiplierStage2Output, flopocoMultiplier232WeightInput, Multiplier232_Output_296);

    MBRightSHR_Float_232_296: entity work.MBRightSHR(rtl)
    GENERIC MAP (96, NumberOfBits)
    PORT MAP (clk, rst, Multiplier232Weight, mbRightSHR232_296Output);

    MB_D_FF_Float_232_296_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR232_296Output, Multiplier232WeightOutput);

    InputIEEE_Float_232_296: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier232WeightOutput, flopocoMultiplier232WeightOutput);

    MB_D_FF_Float_232_296_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier232WeightOutput, flopocoMultiplier232WeightInput);

    MB_D_FF_Float_Multiplier14_236_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier145_Output_181, mb_D_FFMultiplier14_236_0Output);

    MB_D_FF_Float_236_301_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier14_236_0Output, mb_D_FF236_301MultiplierStage1Output);

    MB_D_FF_Float_236_301_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF236_301MultiplierStage1Output, mb_D_FF236_301MultiplierStage2Output);

    Multiplier_Float_236: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF236_301MultiplierStage2Output, flopocoMultiplier236WeightInput, Multiplier236_Output_301);

    MBRightSHR_Float_236_301: entity work.MBRightSHR(rtl)
    GENERIC MAP (89, NumberOfBits)
    PORT MAP (clk, rst, Multiplier236Weight, mbRightSHR236_301Output);

    MB_D_FF_Float_236_301_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR236_301Output, Multiplier236WeightOutput);

    InputIEEE_Float_236_301: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier236WeightOutput, flopocoMultiplier236WeightOutput);

    MB_D_FF_Float_236_301_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier236WeightOutput, flopocoMultiplier236WeightInput);

    MB_D_FF_Float_Multiplier13_237_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier236_Output_301, mb_D_FFMultiplier13_237_0Output);

    MB_D_FF_Float_237_302_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier13_237_0Output, mb_D_FF237_302MultiplierStage1Output);

    MB_D_FF_Float_237_302_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF237_302MultiplierStage1Output, mb_D_FF237_302MultiplierStage2Output);

    Multiplier_Float_237: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF237_302MultiplierStage2Output, flopocoMultiplier237WeightInput, Multiplier237_Output_302);

    MBRightSHR_Float_237_302: entity work.MBRightSHR(rtl)
    GENERIC MAP (96, NumberOfBits)
    PORT MAP (clk, rst, Multiplier237Weight, mbRightSHR237_302Output);

    MB_D_FF_Float_237_302_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR237_302Output, Multiplier237WeightOutput);

    InputIEEE_Float_237_302: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier237WeightOutput, flopocoMultiplier237WeightOutput);

    MB_D_FF_Float_237_302_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier237WeightOutput, flopocoMultiplier237WeightInput);

    MB_D_FF_Float_Adder12_Input1_65_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier237_Output_302, mb_D_FFAdder12_Input1_65_0Output);

    MB_D_FF_Float_65_303_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder12_Input1_65_0Output, mb_D_FF65_303AugendStage1Output);

    MB_D_FF_Float_65_303_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF65_303AugendStage1Output, mb_D_FF65_303AugendStage2Output);

    Adder_Float_65: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF65_303AugendStage2Output, mb_D_FF65_303AddendStage2Output, Adder65_Output_303);

    MB_D_FF_Float_Adder12_Input2_65_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier232_Output_296, mb_D_FFAdder12_Input2_65_0Output);

    MB_D_FF_Float_65_303_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder12_Input2_65_0Output, mb_D_FF65_303AddendStage1Output);

    MB_D_FF_Float_65_303_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF65_303AddendStage1Output, mb_D_FF65_303AddendStage2Output);

    MB_D_FF_Float_Multiplier11_Input1_238_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder65_Output_303, mb_D_FFMultiplier11_Input1_238_0Output);

    MB_D_FF_Float_238_304_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier11_Input1_238_0Output, mb_D_FF238_304MultiplicandStage1Output);

    MB_D_FF_Float_238_304_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF238_304MultiplicandStage1Output, mb_D_FF238_304MultiplicandStage2Output);

    Multiplier_Float_238: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF238_304MultiplicandStage2Output, mb_D_FF238_304MultiplierStage2Output, Multiplier238_Output_304);

    MB_D_FF_Float_Multiplier11_Input2_238_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier227_Output_290, mb_D_FFMultiplier11_Input2_238_0Output);

    MB_D_FF_Float_238_304_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier11_Input2_238_0Output, mb_D_FF238_304MultiplierStage1Output);

    MB_D_FF_Float_238_304_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF238_304MultiplierStage1Output, mb_D_FF238_304MultiplierStage2Output);

    MB_D_FF_Float_Multiplier14_254_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier209_Output_266, mb_D_FFMultiplier14_254_0Output);

    MB_D_FF_Float_254_325_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier14_254_0Output, mb_D_FF254_325MultiplierStage1Output);

    MB_D_FF_Float_254_325_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF254_325MultiplierStage1Output, mb_D_FF254_325MultiplierStage2Output);

    Multiplier_Float_254: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF254_325MultiplierStage2Output, flopocoMultiplier254WeightInput, Multiplier254_Output_325);

    MBRightSHR_Float_254_325: entity work.MBRightSHR(rtl)
    GENERIC MAP (89, NumberOfBits)
    PORT MAP (clk, rst, Multiplier254Weight, mbRightSHR254_325Output);

    MB_D_FF_Float_254_325_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR254_325Output, Multiplier254WeightOutput);

    InputIEEE_Float_254_325: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier254WeightOutput, flopocoMultiplier254WeightOutput);

    MB_D_FF_Float_254_325_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier254WeightOutput, flopocoMultiplier254WeightInput);

    MB_D_FF_Float_Multiplier14_270_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier225_Output_287, mb_D_FFMultiplier14_270_0Output);

    MB_D_FF_Float_270_346_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier14_270_0Output, mb_D_FF270_346MultiplierStage1Output);

    MB_D_FF_Float_270_346_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF270_346MultiplierStage1Output, mb_D_FF270_346MultiplierStage2Output);

    Multiplier_Float_270: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF270_346MultiplierStage2Output, flopocoMultiplier270WeightInput, Multiplier270_Output_346);

    MBRightSHR_Float_270_346: entity work.MBRightSHR(rtl)
    GENERIC MAP (89, NumberOfBits)
    PORT MAP (clk, rst, Multiplier270Weight, mbRightSHR270_346Output);

    MB_D_FF_Float_270_346_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR270_346Output, Multiplier270WeightOutput);

    InputIEEE_Float_270_346: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier270WeightOutput, flopocoMultiplier270WeightOutput);

    MB_D_FF_Float_270_346_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier270WeightOutput, flopocoMultiplier270WeightInput);

    MB_D_FF_Float_Adder13_Input1_76_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier270_Output_346, mb_D_FFAdder13_Input1_76_0Output);

    MB_D_FF_Float_76_347_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder13_Input1_76_0Output, mb_D_FF76_347AugendStage1Output);

    MB_D_FF_Float_76_347_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF76_347AugendStage1Output, mb_D_FF76_347AugendStage2Output);

    Adder_Float_76: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF76_347AugendStage2Output, mb_D_FF76_347AddendStage2Output, Adder76_Output_347);

    MB_D_FF_Float_Adder13_Input2_76_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier254_Output_325, mb_D_FFAdder13_Input2_76_0Output);

    MB_D_FF_Float_76_347_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder13_Input2_76_0Output, mb_D_FF76_347AddendStage1Output);

    MB_D_FF_Float_76_347_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF76_347AddendStage1Output, mb_D_FF76_347AddendStage2Output);

    MB_D_FF_Float_Multiplier12_271_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder76_Output_347, mb_D_FFMultiplier12_271_0Output);

    MB_D_FF_Float_271_348_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier12_271_0Output, mb_D_FF271_348MultiplierStage1Output);

    MB_D_FF_Float_271_348_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF271_348MultiplierStage1Output, mb_D_FF271_348MultiplierStage2Output);

    Multiplier_Float_271: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF271_348MultiplierStage2Output, mb_D_FF271_348MultiplicandStage2Output, Multiplier271_Output_348);

    MBRightSHR_Float_271_348: entity work.MBRightSHR(rtl)
    GENERIC MAP (121, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR271_348Input, mbRightSHR271_348Output);

    MB_D_FF_Float_271_348_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR271_348Output, mb_D_FF271_348MultiplicandStage1Output);

    MB_D_FF_Float_271_348_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF271_348MultiplicandStage1Output, mb_D_FF271_348MultiplicandStage2Output);

    MB_D_FF_Float_Multiplier14_275_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier184_Output_233, mb_D_FFMultiplier14_275_0Output);

    MB_D_FF_Float_275_353_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier14_275_0Output, mb_D_FF275_353MultiplierStage1Output);

    MB_D_FF_Float_275_353_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF275_353MultiplierStage1Output, mb_D_FF275_353MultiplierStage2Output);

    Multiplier_Float_275: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF275_353MultiplierStage2Output, flopocoMultiplier275WeightInput, Multiplier275_Output_353);

    MBRightSHR_Float_275_353: entity work.MBRightSHR(rtl)
    GENERIC MAP (89, NumberOfBits)
    PORT MAP (clk, rst, Multiplier275Weight, mbRightSHR275_353Output);

    MB_D_FF_Float_275_353_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR275_353Output, Multiplier275WeightOutput);

    InputIEEE_Float_275_353: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier275WeightOutput, flopocoMultiplier275WeightOutput);

    MB_D_FF_Float_275_353_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier275WeightOutput, flopocoMultiplier275WeightInput);

    MB_D_FF_Float_Multiplier13_276_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier275_Output_353, mb_D_FFMultiplier13_276_0Output);

    MB_D_FF_Float_276_354_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier13_276_0Output, mb_D_FF276_354MultiplierStage1Output);

    MB_D_FF_Float_276_354_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF276_354MultiplierStage1Output, mb_D_FF276_354MultiplierStage2Output);

    Multiplier_Float_276: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF276_354MultiplierStage2Output, flopocoMultiplier276WeightInput, Multiplier276_Output_354);

    MBRightSHR_Float_276_354: entity work.MBRightSHR(rtl)
    GENERIC MAP (96, NumberOfBits)
    PORT MAP (clk, rst, Multiplier276Weight, mbRightSHR276_354Output);

    MB_D_FF_Float_276_354_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR276_354Output, Multiplier276WeightOutput);

    InputIEEE_Float_276_354: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier276WeightOutput, flopocoMultiplier276WeightOutput);

    MB_D_FF_Float_276_354_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier276WeightOutput, flopocoMultiplier276WeightInput);

    MB_D_FF_Float_Multiplier14_280_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier189_Output_239, mb_D_FFMultiplier14_280_0Output);

    MB_D_FF_Float_280_359_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier14_280_0Output, mb_D_FF280_359MultiplierStage1Output);

    MB_D_FF_Float_280_359_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF280_359MultiplierStage1Output, mb_D_FF280_359MultiplierStage2Output);

    Multiplier_Float_280: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF280_359MultiplierStage2Output, flopocoMultiplier280WeightInput, Multiplier280_Output_359);

    MBRightSHR_Float_280_359: entity work.MBRightSHR(rtl)
    GENERIC MAP (89, NumberOfBits)
    PORT MAP (clk, rst, Multiplier280Weight, mbRightSHR280_359Output);

    MB_D_FF_Float_280_359_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR280_359Output, Multiplier280WeightOutput);

    InputIEEE_Float_280_359: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier280WeightOutput, flopocoMultiplier280WeightOutput);

    MB_D_FF_Float_280_359_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier280WeightOutput, flopocoMultiplier280WeightInput);

    MB_D_FF_Float_Multiplier13_281_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier280_Output_359, mb_D_FFMultiplier13_281_0Output);

    MB_D_FF_Float_281_360_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier13_281_0Output, mb_D_FF281_360MultiplierStage1Output);

    MB_D_FF_Float_281_360_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF281_360MultiplierStage1Output, mb_D_FF281_360MultiplierStage2Output);

    Multiplier_Float_281: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF281_360MultiplierStage2Output, flopocoMultiplier281WeightInput, Multiplier281_Output_360);

    MBRightSHR_Float_281_360: entity work.MBRightSHR(rtl)
    GENERIC MAP (96, NumberOfBits)
    PORT MAP (clk, rst, Multiplier281Weight, mbRightSHR281_360Output);

    MB_D_FF_Float_281_360_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR281_360Output, Multiplier281WeightOutput);

    InputIEEE_Float_281_360: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier281WeightOutput, flopocoMultiplier281WeightOutput);

    MB_D_FF_Float_281_360_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier281WeightOutput, flopocoMultiplier281WeightInput);

    MB_D_FF_Float_Adder12_Input1_79_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier281_Output_360, mb_D_FFAdder12_Input1_79_0Output);

    MB_D_FF_Float_79_361_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder12_Input1_79_0Output, mb_D_FF79_361AugendStage1Output);

    MB_D_FF_Float_79_361_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF79_361AugendStage1Output, mb_D_FF79_361AugendStage2Output);

    Adder_Float_79: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF79_361AugendStage2Output, mb_D_FF79_361AddendStage2Output, Adder79_Output_361);

    MB_D_FF_Float_Adder12_Input2_79_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier276_Output_354, mb_D_FFAdder12_Input2_79_0Output);

    MB_D_FF_Float_79_361_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder12_Input2_79_0Output, mb_D_FF79_361AddendStage1Output);

    MB_D_FF_Float_79_361_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF79_361AddendStage1Output, mb_D_FF79_361AddendStage2Output);

    MB_D_FF_Float_Multiplier11_Input1_282_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder79_Output_361, mb_D_FFMultiplier11_Input1_282_0Output);

    MB_D_FF_Float_282_362_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier11_Input1_282_0Output, mb_D_FF282_362MultiplicandStage1Output);

    MB_D_FF_Float_282_362_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF282_362MultiplicandStage1Output, mb_D_FF282_362MultiplicandStage2Output);

    Multiplier_Float_282: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF282_362MultiplicandStage2Output, mb_D_FF282_362MultiplierStage2Output, Multiplier282_Output_362);

    MB_D_FF_Float_Multiplier11_Input2_282_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier271_Output_348, mb_D_FFMultiplier11_Input2_282_0Output);

    MB_D_FF_Float_282_362_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier11_Input2_282_0Output, mb_D_FF282_362MultiplierStage1Output);

    MB_D_FF_Float_282_362_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF282_362MultiplierStage1Output, mb_D_FF282_362MultiplierStage2Output);

    MB_D_FF_Float_Adder10_Input1_80_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier282_Output_362, mb_D_FFAdder10_Input1_80_0Output);

    MB_D_FF_Float_80_363_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder10_Input1_80_0Output, mb_D_FF80_363AugendStage1Output);

    MB_D_FF_Float_80_363_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF80_363AugendStage1Output, mb_D_FF80_363AugendStage2Output);

    Adder_Float_80: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF80_363AugendStage2Output, mb_D_FF80_363AddendStage2Output, Adder80_Output_363);

    MB_D_FF_Float_Adder10_Input2_80_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier238_Output_304, mb_D_FFAdder10_Input2_80_0Output);

    MB_D_FF_Float_80_363_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder10_Input2_80_0Output, mb_D_FF80_363AddendStage1Output);

    MB_D_FF_Float_80_363_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF80_363AddendStage1Output, mb_D_FF80_363AddendStage2Output);

    MB_D_FF_Float_Multiplier9_283_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder80_Output_363, mb_D_FFMultiplier9_283_0Output);

    MB_D_FF_Float_283_364_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier9_283_0Output, mb_D_FF283_364MultiplierStage1Output);

    MB_D_FF_Float_283_364_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF283_364MultiplierStage1Output, mb_D_FF283_364MultiplierStage2Output);

    Multiplier_Float_283: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF283_364MultiplierStage2Output, mb_D_FF283_364MultiplicandStage2Output, Multiplier283_Output_364);

    MBRightSHR_Float_283_364: entity work.MBRightSHR(rtl)
    GENERIC MAP (160, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR283_364Input, mbRightSHR283_364Output);

    MB_D_FF_Float_283_364_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR283_364Output, mb_D_FF283_364MultiplicandStage1Output);

    MB_D_FF_Float_283_364_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF283_364MultiplicandStage1Output, mb_D_FF283_364MultiplicandStage2Output);

    MB_D_FF_Float_Multiplier8_284_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier283_Output_364, mb_D_FFMultiplier8_284_0Output);

    MB_D_FF_Float_284_365_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier8_284_0Output, mb_D_FF284_365MultiplierStage1Output);

    MB_D_FF_Float_284_365_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF284_365MultiplierStage1Output, mb_D_FF284_365MultiplierStage2Output);

    Multiplier_Float_284: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF284_365MultiplierStage2Output, flopocoMultiplier284WeightInput, Multiplier284_Output_365);

    MBRightSHR_Float_284_365: entity work.MBRightSHR(rtl)
    GENERIC MAP (167, NumberOfBits)
    PORT MAP (clk, rst, Multiplier284Weight, mbRightSHR284_365Output);

    MB_D_FF_Float_284_365_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR284_365Output, Multiplier284WeightOutput);

    InputIEEE_Float_284_365: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier284WeightOutput, flopocoMultiplier284WeightOutput);

    MB_D_FF_Float_284_365_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier284WeightOutput, flopocoMultiplier284WeightInput);

    MB_D_FF_Float_Adder7_Input1_81_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier284_Output_365, mb_D_FFAdder7_Input1_81_0Output);

    MB_D_FF_Float_81_366_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder7_Input1_81_0Output, mb_D_FF81_366AugendStage1Output);

    MB_D_FF_Float_81_366_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF81_366AugendStage1Output, mb_D_FF81_366AugendStage2Output);

    Adder_Float_81: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF81_366AugendStage2Output, mb_D_FF81_366AddendStage2Output, Adder81_Output_366);

    MB_D_FF_Float_Adder7_Input2_81_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier194_Output_246, mb_D_FFAdder7_Input2_81_0Output);

    MB_D_FF_Float_81_366_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder7_Input2_81_0Output, mb_D_FF81_366AddendStage1Output);

    MB_D_FF_Float_81_366_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF81_366AddendStage1Output, mb_D_FF81_366AddendStage2Output);

    MB_D_FF_Float_Multiplier6_Input1_285_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder81_Output_366, mb_D_FFMultiplier6_Input1_285_0Output);

    MB_D_FF_Float_285_367_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier6_Input1_285_0Output, mb_D_FF285_367MultiplicandStage1Output);

    MB_D_FF_Float_285_367_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF285_367MultiplicandStage1Output, mb_D_FF285_367MultiplicandStage2Output);

    Multiplier_Float_285: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF285_367MultiplicandStage2Output, mb_D_FF285_367MultiplierStage2Output, Multiplier285_Output_367);

    MB_D_FF_Float_Multiplier6_Input2_285_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier104_Output_127, mb_D_FFMultiplier6_Input2_285_0Output);

    MB_D_FF_Float_285_367_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier6_Input2_285_0Output, mb_D_FF285_367MultiplierStage1Output);

    MB_D_FF_Float_285_367_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF285_367MultiplierStage1Output, mb_D_FF285_367MultiplierStage2Output);

    MB_D_FF_Float_Multiplier12_310_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier23_Output_28, mb_D_FFMultiplier12_310_0Output);

    MB_D_FF_Float_310_397_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier12_310_0Output, mb_D_FF310_397MultiplierStage1Output);

    MB_D_FF_Float_310_397_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF310_397MultiplierStage1Output, mb_D_FF310_397MultiplierStage2Output);

    Multiplier_Float_310: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF310_397MultiplierStage2Output, flopocoMultiplier310WeightInput, Multiplier310_Output_397);

    MBRightSHR_Float_310_397: entity work.MBRightSHR(rtl)
    GENERIC MAP (121, NumberOfBits)
    PORT MAP (clk, rst, Multiplier310Weight, mbRightSHR310_397Output);

    MB_D_FF_Float_310_397_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR310_397Output, Multiplier310WeightOutput);

    InputIEEE_Float_310_397: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier310WeightOutput, flopocoMultiplier310WeightOutput);

    MB_D_FF_Float_310_397_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier310WeightOutput, flopocoMultiplier310WeightInput);

    MB_D_FF_Float_Multiplier12_335_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier48_Output_58, mb_D_FFMultiplier12_335_0Output);

    MB_D_FF_Float_335_427_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier12_335_0Output, mb_D_FF335_427MultiplierStage1Output);

    MB_D_FF_Float_335_427_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF335_427MultiplierStage1Output, mb_D_FF335_427MultiplierStage2Output);

    Multiplier_Float_335: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF335_427MultiplierStage2Output, flopocoMultiplier335WeightInput, Multiplier335_Output_427);

    MBRightSHR_Float_335_427: entity work.MBRightSHR(rtl)
    GENERIC MAP (121, NumberOfBits)
    PORT MAP (clk, rst, Multiplier335Weight, mbRightSHR335_427Output);

    MB_D_FF_Float_335_427_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR335_427Output, Multiplier335WeightOutput);

    InputIEEE_Float_335_427: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier335WeightOutput, flopocoMultiplier335WeightOutput);

    MB_D_FF_Float_335_427_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier335WeightOutput, flopocoMultiplier335WeightInput);

    MB_D_FF_Float_Adder11_Input1_92_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier335_Output_427, mb_D_FFAdder11_Input1_92_0Output);

    MB_D_FF_Float_92_428_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder11_Input1_92_0Output, mb_D_FF92_428AugendStage1Output);

    MB_D_FF_Float_92_428_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF92_428AugendStage1Output, mb_D_FF92_428AugendStage2Output);

    Adder_Float_92: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF92_428AugendStage2Output, mb_D_FF92_428AddendStage2Output, Adder92_Output_428);

    MB_D_FF_Float_Adder11_Input2_92_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier310_Output_397, mb_D_FFAdder11_Input2_92_0Output);

    MB_D_FF_Float_92_428_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder11_Input2_92_0Output, mb_D_FF92_428AddendStage1Output);

    MB_D_FF_Float_92_428_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF92_428AddendStage1Output, mb_D_FF92_428AddendStage2Output);

    MB_D_FF_Float_Multiplier10_336_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder92_Output_428, mb_D_FFMultiplier10_336_0Output);

    MB_D_FF_Float_336_429_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier10_336_0Output, mb_D_FF336_429MultiplierStage1Output);

    MB_D_FF_Float_336_429_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF336_429MultiplierStage1Output, mb_D_FF336_429MultiplierStage2Output);

    Multiplier_Float_336: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF336_429MultiplierStage2Output, mb_D_FF336_429MultiplicandStage2Output, Multiplier336_Output_429);

    MBRightSHR_Float_336_429: entity work.MBRightSHR(rtl)
    GENERIC MAP (135, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR336_429Input, mbRightSHR336_429Output);

    MB_D_FF_Float_336_429_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR336_429Output, mb_D_FF336_429MultiplicandStage1Output);

    MB_D_FF_Float_336_429_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF336_429MultiplicandStage1Output, mb_D_FF336_429MultiplicandStage2Output);

    MB_D_FF_Float_Multiplier9_337_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier336_Output_429, mb_D_FFMultiplier9_337_0Output);

    MB_D_FF_Float_337_430_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier9_337_0Output, mb_D_FF337_430MultiplierStage1Output);

    MB_D_FF_Float_337_430_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF337_430MultiplierStage1Output, mb_D_FF337_430MultiplierStage2Output);

    Multiplier_Float_337: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF337_430MultiplierStage2Output, flopocoMultiplier337WeightInput, Multiplier337_Output_430);

    MBRightSHR_Float_337_430: entity work.MBRightSHR(rtl)
    GENERIC MAP (160, NumberOfBits)
    PORT MAP (clk, rst, Multiplier337Weight, mbRightSHR337_430Output);

    MB_D_FF_Float_337_430_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR337_430Output, Multiplier337WeightOutput);

    InputIEEE_Float_337_430: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier337WeightOutput, flopocoMultiplier337WeightOutput);

    MB_D_FF_Float_337_430_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier337WeightOutput, flopocoMultiplier337WeightInput);

    MB_D_FF_Float_Multiplier12_362_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier75_Output_91, mb_D_FFMultiplier12_362_0Output);

    MB_D_FF_Float_362_460_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier12_362_0Output, mb_D_FF362_460MultiplierStage1Output);

    MB_D_FF_Float_362_460_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF362_460MultiplierStage1Output, mb_D_FF362_460MultiplierStage2Output);

    Multiplier_Float_362: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF362_460MultiplierStage2Output, flopocoMultiplier362WeightInput, Multiplier362_Output_460);

    MBRightSHR_Float_362_460: entity work.MBRightSHR(rtl)
    GENERIC MAP (121, NumberOfBits)
    PORT MAP (clk, rst, Multiplier362Weight, mbRightSHR362_460Output);

    MB_D_FF_Float_362_460_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR362_460Output, Multiplier362WeightOutput);

    InputIEEE_Float_362_460: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier362WeightOutput, flopocoMultiplier362WeightOutput);

    MB_D_FF_Float_362_460_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier362WeightOutput, flopocoMultiplier362WeightInput);

    MB_D_FF_Float_Multiplier12_387_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier100_Output_121, mb_D_FFMultiplier12_387_0Output);

    MB_D_FF_Float_387_490_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier12_387_0Output, mb_D_FF387_490MultiplierStage1Output);

    MB_D_FF_Float_387_490_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF387_490MultiplierStage1Output, mb_D_FF387_490MultiplierStage2Output);

    Multiplier_Float_387: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF387_490MultiplierStage2Output, flopocoMultiplier387WeightInput, Multiplier387_Output_490);

    MBRightSHR_Float_387_490: entity work.MBRightSHR(rtl)
    GENERIC MAP (121, NumberOfBits)
    PORT MAP (clk, rst, Multiplier387Weight, mbRightSHR387_490Output);

    MB_D_FF_Float_387_490_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR387_490Output, Multiplier387WeightOutput);

    InputIEEE_Float_387_490: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier387WeightOutput, flopocoMultiplier387WeightOutput);

    MB_D_FF_Float_387_490_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier387WeightOutput, flopocoMultiplier387WeightInput);

    MB_D_FF_Float_Adder11_Input1_103_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier387_Output_490, mb_D_FFAdder11_Input1_103_0Output);

    MB_D_FF_Float_103_491_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder11_Input1_103_0Output, mb_D_FF103_491AugendStage1Output);

    MB_D_FF_Float_103_491_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF103_491AugendStage1Output, mb_D_FF103_491AugendStage2Output);

    Adder_Float_103: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF103_491AugendStage2Output, mb_D_FF103_491AddendStage2Output, Adder103_Output_491);

    MB_D_FF_Float_Adder11_Input2_103_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier362_Output_460, mb_D_FFAdder11_Input2_103_0Output);

    MB_D_FF_Float_103_491_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder11_Input2_103_0Output, mb_D_FF103_491AddendStage1Output);

    MB_D_FF_Float_103_491_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF103_491AddendStage1Output, mb_D_FF103_491AddendStage2Output);

    MB_D_FF_Float_Multiplier10_388_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder103_Output_491, mb_D_FFMultiplier10_388_0Output);

    MB_D_FF_Float_388_492_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier10_388_0Output, mb_D_FF388_492MultiplierStage1Output);

    MB_D_FF_Float_388_492_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF388_492MultiplierStage1Output, mb_D_FF388_492MultiplierStage2Output);

    Multiplier_Float_388: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF388_492MultiplierStage2Output, mb_D_FF388_492MultiplicandStage2Output, Multiplier388_Output_492);

    MBRightSHR_Float_388_492: entity work.MBRightSHR(rtl)
    GENERIC MAP (135, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR388_492Input, mbRightSHR388_492Output);

    MB_D_FF_Float_388_492_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR388_492Output, mb_D_FF388_492MultiplicandStage1Output);

    MB_D_FF_Float_388_492_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF388_492MultiplicandStage1Output, mb_D_FF388_492MultiplicandStage2Output);

    MB_D_FF_Float_Multiplier9_389_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier388_Output_492, mb_D_FFMultiplier9_389_0Output);

    MB_D_FF_Float_389_493_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier9_389_0Output, mb_D_FF389_493MultiplierStage1Output);

    MB_D_FF_Float_389_493_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF389_493MultiplierStage1Output, mb_D_FF389_493MultiplierStage2Output);

    Multiplier_Float_389: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF389_493MultiplierStage2Output, flopocoMultiplier389WeightInput, Multiplier389_Output_493);

    MBRightSHR_Float_389_493: entity work.MBRightSHR(rtl)
    GENERIC MAP (160, NumberOfBits)
    PORT MAP (clk, rst, Multiplier389Weight, mbRightSHR389_493Output);

    MB_D_FF_Float_389_493_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR389_493Output, Multiplier389WeightOutput);

    InputIEEE_Float_389_493: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier389WeightOutput, flopocoMultiplier389WeightOutput);

    MB_D_FF_Float_389_493_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier389WeightOutput, flopocoMultiplier389WeightInput);

    MB_D_FF_Float_Adder8_Input1_104_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier389_Output_493, mb_D_FFAdder8_Input1_104_0Output);

    MB_D_FF_Float_104_494_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder8_Input1_104_0Output, mb_D_FF104_494AugendStage1Output);

    MB_D_FF_Float_104_494_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF104_494AugendStage1Output, mb_D_FF104_494AugendStage2Output);

    Adder_Float_104: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF104_494AugendStage2Output, mb_D_FF104_494AddendStage2Output, Adder104_Output_494);

    MB_D_FF_Float_Adder8_Input2_104_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier337_Output_430, mb_D_FFAdder8_Input2_104_0Output);

    MB_D_FF_Float_104_494_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder8_Input2_104_0Output, mb_D_FF104_494AddendStage1Output);

    MB_D_FF_Float_104_494_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF104_494AddendStage1Output, mb_D_FF104_494AddendStage2Output);

    MB_D_FF_Float_Multiplier7_390_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder104_Output_494, mb_D_FFMultiplier7_390_0Output);

    MB_D_FF_Float_390_495_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier7_390_0Output, mb_D_FF390_495MultiplierStage1Output);

    MB_D_FF_Float_390_495_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF390_495MultiplierStage1Output, mb_D_FF390_495MultiplierStage2Output);

    Multiplier_Float_390: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF390_495MultiplierStage2Output, mb_D_FF390_495MultiplicandStage2Output, Multiplier390_Output_495);

    MBRightSHR_Float_390_495: entity work.MBRightSHR(rtl)
    GENERIC MAP (174, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR390_495Input, mbRightSHR390_495Output);

    MB_D_FF_Float_390_495_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR390_495Output, mb_D_FF390_495MultiplicandStage1Output);

    MB_D_FF_Float_390_495_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF390_495MultiplicandStage1Output, mb_D_FF390_495MultiplicandStage2Output);

    MB_D_FF_Float_Multiplier8_480_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier193_Output_245, mb_D_FFMultiplier8_480_0Output);

    MB_D_FF_Float_480_614_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier8_480_0Output, mb_D_FF480_614MultiplierStage1Output);

    MB_D_FF_Float_480_614_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF480_614MultiplierStage1Output, mb_D_FF480_614MultiplierStage2Output);

    Multiplier_Float_480: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF480_614MultiplierStage2Output, flopocoMultiplier480WeightInput, Multiplier480_Output_614);

    MBRightSHR_Float_480_614: entity work.MBRightSHR(rtl)
    GENERIC MAP (167, NumberOfBits)
    PORT MAP (clk, rst, Multiplier480Weight, mbRightSHR480_614Output);

    MB_D_FF_Float_480_614_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR480_614Output, Multiplier480WeightOutput);

    InputIEEE_Float_480_614: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier480WeightOutput, flopocoMultiplier480WeightOutput);

    MB_D_FF_Float_480_614_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier480WeightOutput, flopocoMultiplier480WeightInput);

    MB_D_FF_Float_Multiplier8_570_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier283_Output_364, mb_D_FFMultiplier8_570_0Output);

    MB_D_FF_Float_570_733_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier8_570_0Output, mb_D_FF570_733MultiplierStage1Output);

    MB_D_FF_Float_570_733_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF570_733MultiplierStage1Output, mb_D_FF570_733MultiplierStage2Output);

    Multiplier_Float_570: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF570_733MultiplierStage2Output, flopocoMultiplier570WeightInput, Multiplier570_Output_733);

    MBRightSHR_Float_570_733: entity work.MBRightSHR(rtl)
    GENERIC MAP (167, NumberOfBits)
    PORT MAP (clk, rst, Multiplier570Weight, mbRightSHR570_733Output);

    MB_D_FF_Float_570_733_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR570_733Output, Multiplier570WeightOutput);

    InputIEEE_Float_570_733: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier570WeightOutput, flopocoMultiplier570WeightOutput);

    MB_D_FF_Float_570_733_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier570WeightOutput, flopocoMultiplier570WeightInput);

    MB_D_FF_Float_Adder7_Input1_163_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier570_Output_733, mb_D_FFAdder7_Input1_163_0Output);

    MB_D_FF_Float_163_734_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder7_Input1_163_0Output, mb_D_FF163_734AugendStage1Output);

    MB_D_FF_Float_163_734_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF163_734AugendStage1Output, mb_D_FF163_734AugendStage2Output);

    Adder_Float_163: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF163_734AugendStage2Output, mb_D_FF163_734AddendStage2Output, Adder163_Output_734);

    MB_D_FF_Float_Adder7_Input2_163_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier480_Output_614, mb_D_FFAdder7_Input2_163_0Output);

    MB_D_FF_Float_163_734_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder7_Input2_163_0Output, mb_D_FF163_734AddendStage1Output);

    MB_D_FF_Float_163_734_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF163_734AddendStage1Output, mb_D_FF163_734AddendStage2Output);

    MB_D_FF_Float_Multiplier6_Input1_571_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder163_Output_734, mb_D_FFMultiplier6_Input1_571_0Output);

    MB_D_FF_Float_571_735_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier6_Input1_571_0Output, mb_D_FF571_735MultiplicandStage1Output);

    MB_D_FF_Float_571_735_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF571_735MultiplicandStage1Output, mb_D_FF571_735MultiplicandStage2Output);

    Multiplier_Float_571: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF571_735MultiplicandStage2Output, mb_D_FF571_735MultiplierStage2Output, Multiplier571_Output_735);

    MB_D_FF_Float_Multiplier6_Input2_571_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier390_Output_495, mb_D_FFMultiplier6_Input2_571_0Output);

    MB_D_FF_Float_571_735_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier6_Input2_571_0Output, mb_D_FF571_735MultiplierStage1Output);

    MB_D_FF_Float_571_735_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF571_735MultiplierStage1Output, mb_D_FF571_735MultiplierStage2Output);

    MB_D_FF_Float_Adder5_Input1_164_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier571_Output_735, mb_D_FFAdder5_Input1_164_0Output);

    MB_D_FF_Float_164_736_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder5_Input1_164_0Output, mb_D_FF164_736AugendStage1Output);

    MB_D_FF_Float_164_736_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF164_736AugendStage1Output, mb_D_FF164_736AugendStage2Output);

    Adder_Float_164: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF164_736AugendStage2Output, mb_D_FF164_736AddendStage2Output, Adder164_Output_736);

    MB_D_FF_Float_Adder5_Input2_164_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier285_Output_367, mb_D_FFAdder5_Input2_164_0Output);

    MB_D_FF_Float_164_736_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder5_Input2_164_0Output, mb_D_FF164_736AddendStage1Output);

    MB_D_FF_Float_164_736_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF164_736AddendStage1Output, mb_D_FF164_736AddendStage2Output);

    MB_D_FF_Float_Multiplier4_572_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder164_Output_736, mb_D_FFMultiplier4_572_0Output);

    MB_D_FF_Float_572_737_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier4_572_0Output, mb_D_FF572_737MultiplierStage1Output);

    MB_D_FF_Float_572_737_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF572_737MultiplierStage1Output, mb_D_FF572_737MultiplierStage2Output);

    Multiplier_Float_572: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF572_737MultiplierStage2Output, mb_D_FF572_737MultiplicandStage2Output, Multiplier572_Output_737);

    MBRightSHR_Float_572_737: entity work.MBRightSHR(rtl)
    GENERIC MAP (231, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR572_737Input, mbRightSHR572_737Output);

    MB_D_FF_Float_572_737_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR572_737Output, mb_D_FF572_737MultiplicandStage1Output);

    MB_D_FF_Float_572_737_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF572_737MultiplicandStage1Output, mb_D_FF572_737MultiplicandStage2Output);

    MB_D_FF_Float_Multiplier15_584_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier10_Output_12, mb_D_FFMultiplier15_584_0Output);

    MB_D_FF_Float_584_751_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier15_584_0Output, mb_D_FF584_751MultiplierStage1Output);

    MB_D_FF_Float_584_751_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF584_751MultiplierStage1Output, mb_D_FF584_751MultiplierStage2Output);

    Multiplier_Float_584: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF584_751MultiplierStage2Output, flopocoMultiplier584WeightInput, Multiplier584_Output_751);

    MBRightSHR_Float_584_751: entity work.MBRightSHR(rtl)
    GENERIC MAP (82, NumberOfBits)
    PORT MAP (clk, rst, Multiplier584Weight, mbRightSHR584_751Output);

    MB_D_FF_Float_584_751_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR584_751Output, Multiplier584WeightOutput);

    InputIEEE_Float_584_751: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier584WeightOutput, flopocoMultiplier584WeightOutput);

    MB_D_FF_Float_584_751_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier584WeightOutput, flopocoMultiplier584WeightInput);

    MB_D_FF_Float_Multiplier15_595_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier21_Output_25, mb_D_FFMultiplier15_595_0Output);

    MB_D_FF_Float_595_764_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier15_595_0Output, mb_D_FF595_764MultiplierStage1Output);

    MB_D_FF_Float_595_764_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF595_764MultiplierStage1Output, mb_D_FF595_764MultiplierStage2Output);

    Multiplier_Float_595: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF595_764MultiplierStage2Output, flopocoMultiplier595WeightInput, Multiplier595_Output_764);

    MBRightSHR_Float_595_764: entity work.MBRightSHR(rtl)
    GENERIC MAP (82, NumberOfBits)
    PORT MAP (clk, rst, Multiplier595Weight, mbRightSHR595_764Output);

    MB_D_FF_Float_595_764_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR595_764Output, Multiplier595WeightOutput);

    InputIEEE_Float_595_764: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier595WeightOutput, flopocoMultiplier595WeightOutput);

    MB_D_FF_Float_595_764_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier595WeightOutput, flopocoMultiplier595WeightInput);

    MB_D_FF_Float_Adder14_Input1_169_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier595_Output_764, mb_D_FFAdder14_Input1_169_0Output);

    MB_D_FF_Float_169_765_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder14_Input1_169_0Output, mb_D_FF169_765AugendStage1Output);

    MB_D_FF_Float_169_765_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF169_765AugendStage1Output, mb_D_FF169_765AugendStage2Output);

    Adder_Float_169: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF169_765AugendStage2Output, mb_D_FF169_765AddendStage2Output, Adder169_Output_765);

    MB_D_FF_Float_Adder14_Input2_169_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier584_Output_751, mb_D_FFAdder14_Input2_169_0Output);

    MB_D_FF_Float_169_765_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder14_Input2_169_0Output, mb_D_FF169_765AddendStage1Output);

    MB_D_FF_Float_169_765_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF169_765AddendStage1Output, mb_D_FF169_765AddendStage2Output);

    MB_D_FF_Float_Multiplier13_Input1_596_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder169_Output_765, mb_D_FFMultiplier13_Input1_596_0Output);

    MB_D_FF_Float_596_766_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier13_Input1_596_0Output, mb_D_FF596_766MultiplicandStage1Output);

    MB_D_FF_Float_596_766_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF596_766MultiplicandStage1Output, mb_D_FF596_766MultiplicandStage2Output);

    Multiplier_Float_596: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF596_766MultiplicandStage2Output, mb_D_FF596_766MultiplierStage2Output, Multiplier596_Output_766);

    MB_D_FF_Float_Multiplier13_Input2_596_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier0_Output_0, mb_D_FFMultiplier13_Input2_596_0Output);

    MB_D_FF_Float_596_766_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier13_Input2_596_0Output, mb_D_FF596_766MultiplierStage1Output);

    MB_D_FF_Float_596_766_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF596_766MultiplierStage1Output, mb_D_FF596_766MultiplierStage2Output);

    MB_D_FF_Float_Multiplier12_597_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier596_Output_766, mb_D_FFMultiplier12_597_0Output);

    MB_D_FF_Float_597_767_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier12_597_0Output, mb_D_FF597_767MultiplierStage1Output);

    MB_D_FF_Float_597_767_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF597_767MultiplierStage1Output, mb_D_FF597_767MultiplierStage2Output);

    Multiplier_Float_597: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF597_767MultiplierStage2Output, flopocoMultiplier597WeightInput, Multiplier597_Output_767);

    MBRightSHR_Float_597_767: entity work.MBRightSHR(rtl)
    GENERIC MAP (121, NumberOfBits)
    PORT MAP (clk, rst, Multiplier597Weight, mbRightSHR597_767Output);

    MB_D_FF_Float_597_767_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR597_767Output, Multiplier597WeightOutput);

    InputIEEE_Float_597_767: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier597WeightOutput, flopocoMultiplier597WeightOutput);

    MB_D_FF_Float_597_767_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier597WeightOutput, flopocoMultiplier597WeightInput);

    MB_D_FF_Float_Multiplier15_609_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier35_Output_42, mb_D_FFMultiplier15_609_0Output);

    MB_D_FF_Float_609_781_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier15_609_0Output, mb_D_FF609_781MultiplierStage1Output);

    MB_D_FF_Float_609_781_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF609_781MultiplierStage1Output, mb_D_FF609_781MultiplierStage2Output);

    Multiplier_Float_609: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF609_781MultiplierStage2Output, flopocoMultiplier609WeightInput, Multiplier609_Output_781);

    MBRightSHR_Float_609_781: entity work.MBRightSHR(rtl)
    GENERIC MAP (82, NumberOfBits)
    PORT MAP (clk, rst, Multiplier609Weight, mbRightSHR609_781Output);

    MB_D_FF_Float_609_781_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR609_781Output, Multiplier609WeightOutput);

    InputIEEE_Float_609_781: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier609WeightOutput, flopocoMultiplier609WeightOutput);

    MB_D_FF_Float_609_781_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier609WeightOutput, flopocoMultiplier609WeightInput);

    MB_D_FF_Float_Multiplier15_620_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier46_Output_55, mb_D_FFMultiplier15_620_0Output);

    MB_D_FF_Float_620_794_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier15_620_0Output, mb_D_FF620_794MultiplierStage1Output);

    MB_D_FF_Float_620_794_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF620_794MultiplierStage1Output, mb_D_FF620_794MultiplierStage2Output);

    Multiplier_Float_620: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF620_794MultiplierStage2Output, flopocoMultiplier620WeightInput, Multiplier620_Output_794);

    MBRightSHR_Float_620_794: entity work.MBRightSHR(rtl)
    GENERIC MAP (82, NumberOfBits)
    PORT MAP (clk, rst, Multiplier620Weight, mbRightSHR620_794Output);

    MB_D_FF_Float_620_794_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR620_794Output, Multiplier620WeightOutput);

    InputIEEE_Float_620_794: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier620WeightOutput, flopocoMultiplier620WeightOutput);

    MB_D_FF_Float_620_794_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier620WeightOutput, flopocoMultiplier620WeightInput);

    MB_D_FF_Float_Adder14_Input1_174_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier620_Output_794, mb_D_FFAdder14_Input1_174_0Output);

    MB_D_FF_Float_174_795_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder14_Input1_174_0Output, mb_D_FF174_795AugendStage1Output);

    MB_D_FF_Float_174_795_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF174_795AugendStage1Output, mb_D_FF174_795AugendStage2Output);

    Adder_Float_174: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF174_795AugendStage2Output, mb_D_FF174_795AddendStage2Output, Adder174_Output_795);

    MB_D_FF_Float_Adder14_Input2_174_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier609_Output_781, mb_D_FFAdder14_Input2_174_0Output);

    MB_D_FF_Float_174_795_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder14_Input2_174_0Output, mb_D_FF174_795AddendStage1Output);

    MB_D_FF_Float_174_795_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF174_795AddendStage1Output, mb_D_FF174_795AddendStage2Output);

    MB_D_FF_Float_Multiplier13_Input1_621_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder174_Output_795, mb_D_FFMultiplier13_Input1_621_0Output);

    MB_D_FF_Float_621_796_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier13_Input1_621_0Output, mb_D_FF621_796MultiplicandStage1Output);

    MB_D_FF_Float_621_796_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF621_796MultiplicandStage1Output, mb_D_FF621_796MultiplicandStage2Output);

    Multiplier_Float_621: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF621_796MultiplicandStage2Output, mb_D_FF621_796MultiplierStage2Output, Multiplier621_Output_796);

    MB_D_FF_Float_Multiplier13_Input2_621_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier25_Output_30, mb_D_FFMultiplier13_Input2_621_0Output);

    MB_D_FF_Float_621_796_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier13_Input2_621_0Output, mb_D_FF621_796MultiplierStage1Output);

    MB_D_FF_Float_621_796_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF621_796MultiplierStage1Output, mb_D_FF621_796MultiplierStage2Output);

    MB_D_FF_Float_Multiplier12_622_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier621_Output_796, mb_D_FFMultiplier12_622_0Output);

    MB_D_FF_Float_622_797_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier12_622_0Output, mb_D_FF622_797MultiplierStage1Output);

    MB_D_FF_Float_622_797_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF622_797MultiplierStage1Output, mb_D_FF622_797MultiplierStage2Output);

    Multiplier_Float_622: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF622_797MultiplierStage2Output, flopocoMultiplier622WeightInput, Multiplier622_Output_797);

    MBRightSHR_Float_622_797: entity work.MBRightSHR(rtl)
    GENERIC MAP (121, NumberOfBits)
    PORT MAP (clk, rst, Multiplier622Weight, mbRightSHR622_797Output);

    MB_D_FF_Float_622_797_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR622_797Output, Multiplier622WeightOutput);

    InputIEEE_Float_622_797: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier622WeightOutput, flopocoMultiplier622WeightOutput);

    MB_D_FF_Float_622_797_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier622WeightOutput, flopocoMultiplier622WeightInput);

    MB_D_FF_Float_Adder11_Input1_175_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier622_Output_797, mb_D_FFAdder11_Input1_175_0Output);

    MB_D_FF_Float_175_798_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder11_Input1_175_0Output, mb_D_FF175_798AugendStage1Output);

    MB_D_FF_Float_175_798_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF175_798AugendStage1Output, mb_D_FF175_798AugendStage2Output);

    Adder_Float_175: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF175_798AugendStage2Output, mb_D_FF175_798AddendStage2Output, Adder175_Output_798);

    MB_D_FF_Float_Adder11_Input2_175_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier597_Output_767, mb_D_FFAdder11_Input2_175_0Output);

    MB_D_FF_Float_175_798_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder11_Input2_175_0Output, mb_D_FF175_798AddendStage1Output);

    MB_D_FF_Float_175_798_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF175_798AddendStage1Output, mb_D_FF175_798AddendStage2Output);

    MB_D_FF_Float_Multiplier10_623_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder175_Output_798, mb_D_FFMultiplier10_623_0Output);

    MB_D_FF_Float_623_799_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier10_623_0Output, mb_D_FF623_799MultiplierStage1Output);

    MB_D_FF_Float_623_799_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF623_799MultiplierStage1Output, mb_D_FF623_799MultiplierStage2Output);

    Multiplier_Float_623: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF623_799MultiplierStage2Output, mb_D_FF623_799MultiplicandStage2Output, Multiplier623_Output_799);

    MBRightSHR_Float_623_799: entity work.MBRightSHR(rtl)
    GENERIC MAP (135, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR623_799Input, mbRightSHR623_799Output);

    MB_D_FF_Float_623_799_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR623_799Output, mb_D_FF623_799MultiplicandStage1Output);

    MB_D_FF_Float_623_799_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF623_799MultiplicandStage1Output, mb_D_FF623_799MultiplicandStage2Output);

    MB_D_FF_Float_Multiplier9_624_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier623_Output_799, mb_D_FFMultiplier9_624_0Output);

    MB_D_FF_Float_624_800_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier9_624_0Output, mb_D_FF624_800MultiplierStage1Output);

    MB_D_FF_Float_624_800_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF624_800MultiplierStage1Output, mb_D_FF624_800MultiplierStage2Output);

    Multiplier_Float_624: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF624_800MultiplierStage2Output, flopocoMultiplier624WeightInput, Multiplier624_Output_800);

    MBRightSHR_Float_624_800: entity work.MBRightSHR(rtl)
    GENERIC MAP (160, NumberOfBits)
    PORT MAP (clk, rst, Multiplier624Weight, mbRightSHR624_800Output);

    MB_D_FF_Float_624_800_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR624_800Output, Multiplier624WeightOutput);

    InputIEEE_Float_624_800: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier624WeightOutput, flopocoMultiplier624WeightOutput);

    MB_D_FF_Float_624_800_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier624WeightOutput, flopocoMultiplier624WeightInput);

    MB_D_FF_Float_Multiplier15_636_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier62_Output_75, mb_D_FFMultiplier15_636_0Output);

    MB_D_FF_Float_636_814_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier15_636_0Output, mb_D_FF636_814MultiplierStage1Output);

    MB_D_FF_Float_636_814_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF636_814MultiplierStage1Output, mb_D_FF636_814MultiplierStage2Output);

    Multiplier_Float_636: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF636_814MultiplierStage2Output, flopocoMultiplier636WeightInput, Multiplier636_Output_814);

    MBRightSHR_Float_636_814: entity work.MBRightSHR(rtl)
    GENERIC MAP (82, NumberOfBits)
    PORT MAP (clk, rst, Multiplier636Weight, mbRightSHR636_814Output);

    MB_D_FF_Float_636_814_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR636_814Output, Multiplier636WeightOutput);

    InputIEEE_Float_636_814: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier636WeightOutput, flopocoMultiplier636WeightOutput);

    MB_D_FF_Float_636_814_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier636WeightOutput, flopocoMultiplier636WeightInput);

    MB_D_FF_Float_Multiplier15_647_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier73_Output_88, mb_D_FFMultiplier15_647_0Output);

    MB_D_FF_Float_647_827_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier15_647_0Output, mb_D_FF647_827MultiplierStage1Output);

    MB_D_FF_Float_647_827_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF647_827MultiplierStage1Output, mb_D_FF647_827MultiplierStage2Output);

    Multiplier_Float_647: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF647_827MultiplierStage2Output, flopocoMultiplier647WeightInput, Multiplier647_Output_827);

    MBRightSHR_Float_647_827: entity work.MBRightSHR(rtl)
    GENERIC MAP (82, NumberOfBits)
    PORT MAP (clk, rst, Multiplier647Weight, mbRightSHR647_827Output);

    MB_D_FF_Float_647_827_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR647_827Output, Multiplier647WeightOutput);

    InputIEEE_Float_647_827: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier647WeightOutput, flopocoMultiplier647WeightOutput);

    MB_D_FF_Float_647_827_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier647WeightOutput, flopocoMultiplier647WeightInput);

    MB_D_FF_Float_Adder14_Input1_180_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier647_Output_827, mb_D_FFAdder14_Input1_180_0Output);

    MB_D_FF_Float_180_828_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder14_Input1_180_0Output, mb_D_FF180_828AugendStage1Output);

    MB_D_FF_Float_180_828_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF180_828AugendStage1Output, mb_D_FF180_828AugendStage2Output);

    Adder_Float_180: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF180_828AugendStage2Output, mb_D_FF180_828AddendStage2Output, Adder180_Output_828);

    MB_D_FF_Float_Adder14_Input2_180_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier636_Output_814, mb_D_FFAdder14_Input2_180_0Output);

    MB_D_FF_Float_180_828_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder14_Input2_180_0Output, mb_D_FF180_828AddendStage1Output);

    MB_D_FF_Float_180_828_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF180_828AddendStage1Output, mb_D_FF180_828AddendStage2Output);

    MB_D_FF_Float_Multiplier13_Input1_648_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder180_Output_828, mb_D_FFMultiplier13_Input1_648_0Output);

    MB_D_FF_Float_648_829_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier13_Input1_648_0Output, mb_D_FF648_829MultiplicandStage1Output);

    MB_D_FF_Float_648_829_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF648_829MultiplicandStage1Output, mb_D_FF648_829MultiplicandStage2Output);

    Multiplier_Float_648: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF648_829MultiplicandStage2Output, mb_D_FF648_829MultiplierStage2Output, Multiplier648_Output_829);

    MB_D_FF_Float_Multiplier13_Input2_648_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier0_Output_0, mb_D_FFMultiplier13_Input2_648_0Output);

    MB_D_FF_Float_648_829_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier13_Input2_648_0Output, mb_D_FF648_829MultiplierStage1Output);

    MB_D_FF_Float_648_829_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF648_829MultiplierStage1Output, mb_D_FF648_829MultiplierStage2Output);

    MB_D_FF_Float_Multiplier12_649_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier648_Output_829, mb_D_FFMultiplier12_649_0Output);

    MB_D_FF_Float_649_830_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier12_649_0Output, mb_D_FF649_830MultiplierStage1Output);

    MB_D_FF_Float_649_830_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF649_830MultiplierStage1Output, mb_D_FF649_830MultiplierStage2Output);

    Multiplier_Float_649: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF649_830MultiplierStage2Output, flopocoMultiplier649WeightInput, Multiplier649_Output_830);

    MBRightSHR_Float_649_830: entity work.MBRightSHR(rtl)
    GENERIC MAP (121, NumberOfBits)
    PORT MAP (clk, rst, Multiplier649Weight, mbRightSHR649_830Output);

    MB_D_FF_Float_649_830_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR649_830Output, Multiplier649WeightOutput);

    InputIEEE_Float_649_830: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier649WeightOutput, flopocoMultiplier649WeightOutput);

    MB_D_FF_Float_649_830_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier649WeightOutput, flopocoMultiplier649WeightInput);

    MB_D_FF_Float_Multiplier15_661_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier87_Output_105, mb_D_FFMultiplier15_661_0Output);

    MB_D_FF_Float_661_844_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier15_661_0Output, mb_D_FF661_844MultiplierStage1Output);

    MB_D_FF_Float_661_844_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF661_844MultiplierStage1Output, mb_D_FF661_844MultiplierStage2Output);

    Multiplier_Float_661: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF661_844MultiplierStage2Output, flopocoMultiplier661WeightInput, Multiplier661_Output_844);

    MBRightSHR_Float_661_844: entity work.MBRightSHR(rtl)
    GENERIC MAP (82, NumberOfBits)
    PORT MAP (clk, rst, Multiplier661Weight, mbRightSHR661_844Output);

    MB_D_FF_Float_661_844_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR661_844Output, Multiplier661WeightOutput);

    InputIEEE_Float_661_844: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier661WeightOutput, flopocoMultiplier661WeightOutput);

    MB_D_FF_Float_661_844_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier661WeightOutput, flopocoMultiplier661WeightInput);

    MB_D_FF_Float_Multiplier15_672_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier98_Output_118, mb_D_FFMultiplier15_672_0Output);

    MB_D_FF_Float_672_857_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier15_672_0Output, mb_D_FF672_857MultiplierStage1Output);

    MB_D_FF_Float_672_857_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF672_857MultiplierStage1Output, mb_D_FF672_857MultiplierStage2Output);

    Multiplier_Float_672: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF672_857MultiplierStage2Output, flopocoMultiplier672WeightInput, Multiplier672_Output_857);

    MBRightSHR_Float_672_857: entity work.MBRightSHR(rtl)
    GENERIC MAP (82, NumberOfBits)
    PORT MAP (clk, rst, Multiplier672Weight, mbRightSHR672_857Output);

    MB_D_FF_Float_672_857_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR672_857Output, Multiplier672WeightOutput);

    InputIEEE_Float_672_857: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier672WeightOutput, flopocoMultiplier672WeightOutput);

    MB_D_FF_Float_672_857_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier672WeightOutput, flopocoMultiplier672WeightInput);

    MB_D_FF_Float_Adder14_Input1_185_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier672_Output_857, mb_D_FFAdder14_Input1_185_0Output);

    MB_D_FF_Float_185_858_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder14_Input1_185_0Output, mb_D_FF185_858AugendStage1Output);

    MB_D_FF_Float_185_858_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF185_858AugendStage1Output, mb_D_FF185_858AugendStage2Output);

    Adder_Float_185: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF185_858AugendStage2Output, mb_D_FF185_858AddendStage2Output, Adder185_Output_858);

    MB_D_FF_Float_Adder14_Input2_185_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier661_Output_844, mb_D_FFAdder14_Input2_185_0Output);

    MB_D_FF_Float_185_858_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder14_Input2_185_0Output, mb_D_FF185_858AddendStage1Output);

    MB_D_FF_Float_185_858_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF185_858AddendStage1Output, mb_D_FF185_858AddendStage2Output);

    MB_D_FF_Float_Multiplier13_Input1_673_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder185_Output_858, mb_D_FFMultiplier13_Input1_673_0Output);

    MB_D_FF_Float_673_859_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier13_Input1_673_0Output, mb_D_FF673_859MultiplicandStage1Output);

    MB_D_FF_Float_673_859_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF673_859MultiplicandStage1Output, mb_D_FF673_859MultiplicandStage2Output);

    Multiplier_Float_673: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF673_859MultiplicandStage2Output, mb_D_FF673_859MultiplierStage2Output, Multiplier673_Output_859);

    MB_D_FF_Float_Multiplier13_Input2_673_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier25_Output_30, mb_D_FFMultiplier13_Input2_673_0Output);

    MB_D_FF_Float_673_859_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier13_Input2_673_0Output, mb_D_FF673_859MultiplierStage1Output);

    MB_D_FF_Float_673_859_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF673_859MultiplierStage1Output, mb_D_FF673_859MultiplierStage2Output);

    MB_D_FF_Float_Multiplier12_674_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier673_Output_859, mb_D_FFMultiplier12_674_0Output);

    MB_D_FF_Float_674_860_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier12_674_0Output, mb_D_FF674_860MultiplierStage1Output);

    MB_D_FF_Float_674_860_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF674_860MultiplierStage1Output, mb_D_FF674_860MultiplierStage2Output);

    Multiplier_Float_674: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF674_860MultiplierStage2Output, flopocoMultiplier674WeightInput, Multiplier674_Output_860);

    MBRightSHR_Float_674_860: entity work.MBRightSHR(rtl)
    GENERIC MAP (121, NumberOfBits)
    PORT MAP (clk, rst, Multiplier674Weight, mbRightSHR674_860Output);

    MB_D_FF_Float_674_860_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR674_860Output, Multiplier674WeightOutput);

    InputIEEE_Float_674_860: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier674WeightOutput, flopocoMultiplier674WeightOutput);

    MB_D_FF_Float_674_860_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier674WeightOutput, flopocoMultiplier674WeightInput);

    MB_D_FF_Float_Adder11_Input1_186_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier674_Output_860, mb_D_FFAdder11_Input1_186_0Output);

    MB_D_FF_Float_186_861_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder11_Input1_186_0Output, mb_D_FF186_861AugendStage1Output);

    MB_D_FF_Float_186_861_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF186_861AugendStage1Output, mb_D_FF186_861AugendStage2Output);

    Adder_Float_186: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF186_861AugendStage2Output, mb_D_FF186_861AddendStage2Output, Adder186_Output_861);

    MB_D_FF_Float_Adder11_Input2_186_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier649_Output_830, mb_D_FFAdder11_Input2_186_0Output);

    MB_D_FF_Float_186_861_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder11_Input2_186_0Output, mb_D_FF186_861AddendStage1Output);

    MB_D_FF_Float_186_861_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF186_861AddendStage1Output, mb_D_FF186_861AddendStage2Output);

    MB_D_FF_Float_Multiplier10_675_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder186_Output_861, mb_D_FFMultiplier10_675_0Output);

    MB_D_FF_Float_675_862_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier10_675_0Output, mb_D_FF675_862MultiplierStage1Output);

    MB_D_FF_Float_675_862_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF675_862MultiplierStage1Output, mb_D_FF675_862MultiplierStage2Output);

    Multiplier_Float_675: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF675_862MultiplierStage2Output, mb_D_FF675_862MultiplicandStage2Output, Multiplier675_Output_862);

    MBRightSHR_Float_675_862: entity work.MBRightSHR(rtl)
    GENERIC MAP (135, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR675_862Input, mbRightSHR675_862Output);

    MB_D_FF_Float_675_862_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR675_862Output, mb_D_FF675_862MultiplicandStage1Output);

    MB_D_FF_Float_675_862_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF675_862MultiplicandStage1Output, mb_D_FF675_862MultiplicandStage2Output);

    MB_D_FF_Float_Multiplier9_676_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier675_Output_862, mb_D_FFMultiplier9_676_0Output);

    MB_D_FF_Float_676_863_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier9_676_0Output, mb_D_FF676_863MultiplierStage1Output);

    MB_D_FF_Float_676_863_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF676_863MultiplierStage1Output, mb_D_FF676_863MultiplierStage2Output);

    Multiplier_Float_676: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF676_863MultiplierStage2Output, flopocoMultiplier676WeightInput, Multiplier676_Output_863);

    MBRightSHR_Float_676_863: entity work.MBRightSHR(rtl)
    GENERIC MAP (160, NumberOfBits)
    PORT MAP (clk, rst, Multiplier676Weight, mbRightSHR676_863Output);

    MB_D_FF_Float_676_863_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR676_863Output, Multiplier676WeightOutput);

    InputIEEE_Float_676_863: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier676WeightOutput, flopocoMultiplier676WeightOutput);

    MB_D_FF_Float_676_863_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier676WeightOutput, flopocoMultiplier676WeightInput);

    MB_D_FF_Float_Adder8_Input1_187_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier676_Output_863, mb_D_FFAdder8_Input1_187_0Output);

    MB_D_FF_Float_187_864_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder8_Input1_187_0Output, mb_D_FF187_864AugendStage1Output);

    MB_D_FF_Float_187_864_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF187_864AugendStage1Output, mb_D_FF187_864AugendStage2Output);

    Adder_Float_187: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF187_864AugendStage2Output, mb_D_FF187_864AddendStage2Output, Adder187_Output_864);

    MB_D_FF_Float_Adder8_Input2_187_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier624_Output_800, mb_D_FFAdder8_Input2_187_0Output);

    MB_D_FF_Float_187_864_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder8_Input2_187_0Output, mb_D_FF187_864AddendStage1Output);

    MB_D_FF_Float_187_864_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF187_864AddendStage1Output, mb_D_FF187_864AddendStage2Output);

    MB_D_FF_Float_Multiplier7_677_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder187_Output_864, mb_D_FFMultiplier7_677_0Output);

    MB_D_FF_Float_677_865_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier7_677_0Output, mb_D_FF677_865MultiplierStage1Output);

    MB_D_FF_Float_677_865_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF677_865MultiplierStage1Output, mb_D_FF677_865MultiplierStage2Output);

    Multiplier_Float_677: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF677_865MultiplierStage2Output, mb_D_FF677_865MultiplicandStage2Output, Multiplier677_Output_865);

    MBRightSHR_Float_677_865: entity work.MBRightSHR(rtl)
    GENERIC MAP (174, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR677_865Input, mbRightSHR677_865Output);

    MB_D_FF_Float_677_865_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR677_865Output, mb_D_FF677_865MultiplicandStage1Output);

    MB_D_FF_Float_677_865_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF677_865MultiplicandStage1Output, mb_D_FF677_865MultiplicandStage2Output);

    MBRightSHR_Float_678_866: entity work.MBRightSHR(rtl)
    GENERIC MAP (4, NumberOfBits)
    PORT MAP (clk, rst, Multiplier678Weight, mbRightSHR678_866Output);

    MB_D_FF_Float_678_866_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR678_866Output, Multiplier678WeightOutput);

    InputIEEE_Float_678_866: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier678WeightOutput, flopocoMultiplier678WeightOutput);

    MB_D_FF_Float_678_866_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier678WeightOutput, flopocoMultiplier678WeightInput);

    Multiplier_Float_678: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier678WeightInput, mb_D_FF678_866MultiplierStage2Output, Multiplier678_Output_866);

    MB_D_FF_Float_Multiplier21_678_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier21_678_0Input, mb_D_FFMultiplier21_678_0Output);

    MB_D_FF_Float_678_866_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier21_678_0Output, mb_D_FF678_866MultiplierStage1Output);

    MB_D_FF_Float_678_866_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF678_866MultiplierStage1Output, mb_D_FF678_866MultiplierStage2Output);

    MBRightSHR_Float_679_867: entity work.MBRightSHR(rtl)
    GENERIC MAP (4, NumberOfBits)
    PORT MAP (clk, rst, Multiplier679Weight, mbRightSHR679_867Output);

    MB_D_FF_Float_679_867_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR679_867Output, Multiplier679WeightOutput);

    InputIEEE_Float_679_867: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier679WeightOutput, flopocoMultiplier679WeightOutput);

    MB_D_FF_Float_679_867_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier679WeightOutput, flopocoMultiplier679WeightInput);

    Multiplier_Float_679: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier679WeightInput, mb_D_FF679_867MultiplierStage2Output, Multiplier679_Output_867);

    MB_D_FF_Float_Multiplier21_679_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier21_679_0Input, mb_D_FFMultiplier21_679_0Output);

    MB_D_FF_Float_679_867_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier21_679_0Output, mb_D_FF679_867MultiplierStage1Output);

    MB_D_FF_Float_679_867_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF679_867MultiplierStage1Output, mb_D_FF679_867MultiplierStage2Output);

    MB_D_FF_Float_Adder20_Input1_188_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier679_Output_867, mb_D_FFAdder20_Input1_188_0Output);

    MB_D_FF_Float_188_868_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder20_Input1_188_0Output, mb_D_FF188_868AugendStage1Output);

    MB_D_FF_Float_188_868_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF188_868AugendStage1Output, mb_D_FF188_868AugendStage2Output);

    Adder_Float_188: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF188_868AugendStage2Output, mb_D_FF188_868AddendStage2Output, Adder188_Output_868);

    MB_D_FF_Float_Adder20_Input2_188_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier678_Output_866, mb_D_FFAdder20_Input2_188_0Output);

    MB_D_FF_Float_188_868_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder20_Input2_188_0Output, mb_D_FF188_868AddendStage1Output);

    MB_D_FF_Float_188_868_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF188_868AddendStage1Output, mb_D_FF188_868AddendStage2Output);

    MB_D_FF_Float_Multiplier19_680_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder188_Output_868, mb_D_FFMultiplier19_680_0Output);

    MB_D_FF_Float_680_869_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier19_680_0Output, mb_D_FF680_869MultiplierStage1Output);

    MB_D_FF_Float_680_869_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF680_869MultiplierStage1Output, mb_D_FF680_869MultiplierStage2Output);

    Multiplier_Float_680: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF680_869MultiplierStage2Output, mb_D_FF680_869MultiplicandStage2Output, Multiplier680_Output_869);

    MBRightSHR_Float_680_869: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR680_869Input, mbRightSHR680_869Output);

    MB_D_FF_Float_680_869_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR680_869Output, mb_D_FF680_869MultiplicandStage1Output);

    MB_D_FF_Float_680_869_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF680_869MultiplicandStage1Output, mb_D_FF680_869MultiplicandStage2Output);

    MB_D_FF_Float_Multiplier18_681_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier680_Output_869, mb_D_FFMultiplier18_681_0Output);

    MB_D_FF_Float_681_870_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier18_681_0Output, mb_D_FF681_870MultiplierStage1Output);

    MB_D_FF_Float_681_870_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF681_870MultiplierStage1Output, mb_D_FF681_870MultiplierStage2Output);

    Multiplier_Float_681: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF681_870MultiplierStage2Output, flopocoMultiplier681WeightInput, Multiplier681_Output_870);

    MBRightSHR_Float_681_870: entity work.MBRightSHR(rtl)
    GENERIC MAP (43, NumberOfBits)
    PORT MAP (clk, rst, Multiplier681Weight, mbRightSHR681_870Output);

    MB_D_FF_Float_681_870_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR681_870Output, Multiplier681WeightOutput);

    InputIEEE_Float_681_870: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier681WeightOutput, flopocoMultiplier681WeightOutput);

    MB_D_FF_Float_681_870_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier681WeightOutput, flopocoMultiplier681WeightInput);

    MB_D_FF_Float_Multiplier17_Input1_684_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder24_Output_135, mb_D_FFMultiplier17_Input1_684_0Output);

    MB_D_FF_Float_684_874_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier17_Input1_684_0Output, mb_D_FF684_874MultiplicandStage1Output);

    MB_D_FF_Float_684_874_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF684_874MultiplicandStage1Output, mb_D_FF684_874MultiplicandStage2Output);

    Multiplier_Float_684: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF684_874MultiplicandStage2Output, mb_D_FF684_874MultiplierStage2Output, Multiplier684_Output_874);

    MB_D_FF_Float_Multiplier17_Input2_684_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier681_Output_870, mb_D_FFMultiplier17_Input2_684_0Output);

    MB_D_FF_Float_684_874_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier17_Input2_684_0Output, mb_D_FF684_874MultiplierStage1Output);

    MB_D_FF_Float_684_874_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF684_874MultiplierStage1Output, mb_D_FF684_874MultiplierStage2Output);

    MBRightSHR_Float_685_875: entity work.MBRightSHR(rtl)
    GENERIC MAP (4, NumberOfBits)
    PORT MAP (clk, rst, Multiplier685Weight, mbRightSHR685_875Output);

    MB_D_FF_Float_685_875_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR685_875Output, Multiplier685WeightOutput);

    InputIEEE_Float_685_875: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier685WeightOutput, flopocoMultiplier685WeightOutput);

    MB_D_FF_Float_685_875_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier685WeightOutput, flopocoMultiplier685WeightInput);

    Multiplier_Float_685: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier685WeightInput, mb_D_FF685_875MultiplierStage2Output, Multiplier685_Output_875);

    MB_D_FF_Float_Multiplier21_685_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier21_685_0Input, mb_D_FFMultiplier21_685_0Output);

    MB_D_FF_Float_685_875_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier21_685_0Output, mb_D_FF685_875MultiplierStage1Output);

    MB_D_FF_Float_685_875_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF685_875MultiplierStage1Output, mb_D_FF685_875MultiplierStage2Output);

    MBRightSHR_Float_686_876: entity work.MBRightSHR(rtl)
    GENERIC MAP (4, NumberOfBits)
    PORT MAP (clk, rst, Multiplier686Weight, mbRightSHR686_876Output);

    MB_D_FF_Float_686_876_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR686_876Output, Multiplier686WeightOutput);

    InputIEEE_Float_686_876: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier686WeightOutput, flopocoMultiplier686WeightOutput);

    MB_D_FF_Float_686_876_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier686WeightOutput, flopocoMultiplier686WeightInput);

    Multiplier_Float_686: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier686WeightInput, mb_D_FF686_876MultiplierStage2Output, Multiplier686_Output_876);

    MB_D_FF_Float_Multiplier21_686_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier21_686_0Input, mb_D_FFMultiplier21_686_0Output);

    MB_D_FF_Float_686_876_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier21_686_0Output, mb_D_FF686_876MultiplierStage1Output);

    MB_D_FF_Float_686_876_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF686_876MultiplierStage1Output, mb_D_FF686_876MultiplierStage2Output);

    MB_D_FF_Float_Adder20_Input1_190_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier686_Output_876, mb_D_FFAdder20_Input1_190_0Output);

    MB_D_FF_Float_190_877_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder20_Input1_190_0Output, mb_D_FF190_877AugendStage1Output);

    MB_D_FF_Float_190_877_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF190_877AugendStage1Output, mb_D_FF190_877AugendStage2Output);

    Adder_Float_190: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF190_877AugendStage2Output, mb_D_FF190_877AddendStage2Output, Adder190_Output_877);

    MB_D_FF_Float_Adder20_Input2_190_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier685_Output_875, mb_D_FFAdder20_Input2_190_0Output);

    MB_D_FF_Float_190_877_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder20_Input2_190_0Output, mb_D_FF190_877AddendStage1Output);

    MB_D_FF_Float_190_877_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF190_877AddendStage1Output, mb_D_FF190_877AddendStage2Output);

    MB_D_FF_Float_Multiplier19_687_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder190_Output_877, mb_D_FFMultiplier19_687_0Output);

    MB_D_FF_Float_687_878_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier19_687_0Output, mb_D_FF687_878MultiplierStage1Output);

    MB_D_FF_Float_687_878_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF687_878MultiplierStage1Output, mb_D_FF687_878MultiplierStage2Output);

    Multiplier_Float_687: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF687_878MultiplierStage2Output, mb_D_FF687_878MultiplicandStage2Output, Multiplier687_Output_878);

    MBRightSHR_Float_687_878: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR687_878Input, mbRightSHR687_878Output);

    MB_D_FF_Float_687_878_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR687_878Output, mb_D_FF687_878MultiplicandStage1Output);

    MB_D_FF_Float_687_878_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF687_878MultiplicandStage1Output, mb_D_FF687_878MultiplicandStage2Output);

    MB_D_FF_Float_Multiplier18_688_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier687_Output_878, mb_D_FFMultiplier18_688_0Output);

    MB_D_FF_Float_688_879_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier18_688_0Output, mb_D_FF688_879MultiplierStage1Output);

    MB_D_FF_Float_688_879_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF688_879MultiplierStage1Output, mb_D_FF688_879MultiplierStage2Output);

    Multiplier_Float_688: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF688_879MultiplierStage2Output, flopocoMultiplier688WeightInput, Multiplier688_Output_879);

    MBRightSHR_Float_688_879: entity work.MBRightSHR(rtl)
    GENERIC MAP (43, NumberOfBits)
    PORT MAP (clk, rst, Multiplier688Weight, mbRightSHR688_879Output);

    MB_D_FF_Float_688_879_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR688_879Output, Multiplier688WeightOutput);

    InputIEEE_Float_688_879: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier688WeightOutput, flopocoMultiplier688WeightOutput);

    MB_D_FF_Float_688_879_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier688WeightOutput, flopocoMultiplier688WeightInput);

    MB_D_FF_Float_Multiplier17_Input1_691_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder26_Output_144, mb_D_FFMultiplier17_Input1_691_0Output);

    MB_D_FF_Float_691_883_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier17_Input1_691_0Output, mb_D_FF691_883MultiplicandStage1Output);

    MB_D_FF_Float_691_883_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF691_883MultiplicandStage1Output, mb_D_FF691_883MultiplicandStage2Output);

    Multiplier_Float_691: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF691_883MultiplicandStage2Output, mb_D_FF691_883MultiplierStage2Output, Multiplier691_Output_883);

    MB_D_FF_Float_Multiplier17_Input2_691_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier688_Output_879, mb_D_FFMultiplier17_Input2_691_0Output);

    MB_D_FF_Float_691_883_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier17_Input2_691_0Output, mb_D_FF691_883MultiplierStage1Output);

    MB_D_FF_Float_691_883_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF691_883MultiplierStage1Output, mb_D_FF691_883MultiplierStage2Output);

    MB_D_FF_Float_Adder16_Input1_192_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier691_Output_883, mb_D_FFAdder16_Input1_192_0Output);

    MB_D_FF_Float_192_884_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder16_Input1_192_0Output, mb_D_FF192_884AugendStage1Output);

    MB_D_FF_Float_192_884_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF192_884AugendStage1Output, mb_D_FF192_884AugendStage2Output);

    Adder_Float_192: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF192_884AugendStage2Output, mb_D_FF192_884AddendStage2Output, Adder192_Output_884);

    MB_D_FF_Float_Adder16_Input2_192_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier684_Output_874, mb_D_FFAdder16_Input2_192_0Output);

    MB_D_FF_Float_192_884_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder16_Input2_192_0Output, mb_D_FF192_884AddendStage1Output);

    MB_D_FF_Float_192_884_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF192_884AddendStage1Output, mb_D_FF192_884AddendStage2Output);

    MB_D_FF_Float_Multiplier15_692_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder192_Output_884, mb_D_FFMultiplier15_692_0Output);

    MB_D_FF_Float_692_885_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier15_692_0Output, mb_D_FF692_885MultiplierStage1Output);

    MB_D_FF_Float_692_885_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF692_885MultiplierStage1Output, mb_D_FF692_885MultiplierStage2Output);

    Multiplier_Float_692: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF692_885MultiplierStage2Output, mb_D_FF692_885MultiplicandStage2Output, Multiplier692_Output_885);

    MBRightSHR_Float_692_885: entity work.MBRightSHR(rtl)
    GENERIC MAP (82, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR692_885Input, mbRightSHR692_885Output);

    MB_D_FF_Float_692_885_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR692_885Output, mb_D_FF692_885MultiplicandStage1Output);

    MB_D_FF_Float_692_885_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF692_885MultiplicandStage1Output, mb_D_FF692_885MultiplicandStage2Output);

    MB_D_FF_Float_Multiplier14_693_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier692_Output_885, mb_D_FFMultiplier14_693_0Output);

    MB_D_FF_Float_693_886_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier14_693_0Output, mb_D_FF693_886MultiplierStage1Output);

    MB_D_FF_Float_693_886_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF693_886MultiplierStage1Output, mb_D_FF693_886MultiplierStage2Output);

    Multiplier_Float_693: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF693_886MultiplierStage2Output, flopocoMultiplier693WeightInput, Multiplier693_Output_886);

    MBRightSHR_Float_693_886: entity work.MBRightSHR(rtl)
    GENERIC MAP (89, NumberOfBits)
    PORT MAP (clk, rst, Multiplier693Weight, mbRightSHR693_886Output);

    MB_D_FF_Float_693_886_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR693_886Output, Multiplier693WeightOutput);

    InputIEEE_Float_693_886: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier693WeightOutput, flopocoMultiplier693WeightOutput);

    MB_D_FF_Float_693_886_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier693WeightOutput, flopocoMultiplier693WeightInput);

    MBRightSHR_Float_694_887: entity work.MBRightSHR(rtl)
    GENERIC MAP (4, NumberOfBits)
    PORT MAP (clk, rst, Multiplier694Weight, mbRightSHR694_887Output);

    MB_D_FF_Float_694_887_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR694_887Output, Multiplier694WeightOutput);

    InputIEEE_Float_694_887: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier694WeightOutput, flopocoMultiplier694WeightOutput);

    MB_D_FF_Float_694_887_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier694WeightOutput, flopocoMultiplier694WeightInput);

    Multiplier_Float_694: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier694WeightInput, mb_D_FF694_887MultiplierStage2Output, Multiplier694_Output_887);

    MB_D_FF_Float_Multiplier21_694_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier21_694_0Input, mb_D_FFMultiplier21_694_0Output);

    MB_D_FF_Float_694_887_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier21_694_0Output, mb_D_FF694_887MultiplierStage1Output);

    MB_D_FF_Float_694_887_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF694_887MultiplierStage1Output, mb_D_FF694_887MultiplierStage2Output);

    MBRightSHR_Float_695_888: entity work.MBRightSHR(rtl)
    GENERIC MAP (4, NumberOfBits)
    PORT MAP (clk, rst, Multiplier695Weight, mbRightSHR695_888Output);

    MB_D_FF_Float_695_888_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR695_888Output, Multiplier695WeightOutput);

    InputIEEE_Float_695_888: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier695WeightOutput, flopocoMultiplier695WeightOutput);

    MB_D_FF_Float_695_888_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier695WeightOutput, flopocoMultiplier695WeightInput);

    Multiplier_Float_695: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier695WeightInput, mb_D_FF695_888MultiplierStage2Output, Multiplier695_Output_888);

    MB_D_FF_Float_Multiplier21_695_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier21_695_0Input, mb_D_FFMultiplier21_695_0Output);

    MB_D_FF_Float_695_888_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier21_695_0Output, mb_D_FF695_888MultiplierStage1Output);

    MB_D_FF_Float_695_888_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF695_888MultiplierStage1Output, mb_D_FF695_888MultiplierStage2Output);

    MB_D_FF_Float_Adder20_Input1_193_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier695_Output_888, mb_D_FFAdder20_Input1_193_0Output);

    MB_D_FF_Float_193_889_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder20_Input1_193_0Output, mb_D_FF193_889AugendStage1Output);

    MB_D_FF_Float_193_889_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF193_889AugendStage1Output, mb_D_FF193_889AugendStage2Output);

    Adder_Float_193: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF193_889AugendStage2Output, mb_D_FF193_889AddendStage2Output, Adder193_Output_889);

    MB_D_FF_Float_Adder20_Input2_193_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier694_Output_887, mb_D_FFAdder20_Input2_193_0Output);

    MB_D_FF_Float_193_889_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder20_Input2_193_0Output, mb_D_FF193_889AddendStage1Output);

    MB_D_FF_Float_193_889_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF193_889AddendStage1Output, mb_D_FF193_889AddendStage2Output);

    MB_D_FF_Float_Multiplier19_696_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder193_Output_889, mb_D_FFMultiplier19_696_0Output);

    MB_D_FF_Float_696_890_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier19_696_0Output, mb_D_FF696_890MultiplierStage1Output);

    MB_D_FF_Float_696_890_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF696_890MultiplierStage1Output, mb_D_FF696_890MultiplierStage2Output);

    Multiplier_Float_696: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF696_890MultiplierStage2Output, mb_D_FF696_890MultiplicandStage2Output, Multiplier696_Output_890);

    MBRightSHR_Float_696_890: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR696_890Input, mbRightSHR696_890Output);

    MB_D_FF_Float_696_890_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR696_890Output, mb_D_FF696_890MultiplicandStage1Output);

    MB_D_FF_Float_696_890_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF696_890MultiplicandStage1Output, mb_D_FF696_890MultiplicandStage2Output);

    MB_D_FF_Float_Multiplier18_697_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier696_Output_890, mb_D_FFMultiplier18_697_0Output);

    MB_D_FF_Float_697_891_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier18_697_0Output, mb_D_FF697_891MultiplierStage1Output);

    MB_D_FF_Float_697_891_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF697_891MultiplierStage1Output, mb_D_FF697_891MultiplierStage2Output);

    Multiplier_Float_697: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF697_891MultiplierStage2Output, flopocoMultiplier697WeightInput, Multiplier697_Output_891);

    MBRightSHR_Float_697_891: entity work.MBRightSHR(rtl)
    GENERIC MAP (43, NumberOfBits)
    PORT MAP (clk, rst, Multiplier697Weight, mbRightSHR697_891Output);

    MB_D_FF_Float_697_891_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR697_891Output, Multiplier697WeightOutput);

    InputIEEE_Float_697_891: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier697WeightOutput, flopocoMultiplier697WeightOutput);

    MB_D_FF_Float_697_891_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier697WeightOutput, flopocoMultiplier697WeightInput);

    MB_D_FF_Float_Multiplier17_Input1_700_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder29_Output_156, mb_D_FFMultiplier17_Input1_700_0Output);

    MB_D_FF_Float_700_895_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier17_Input1_700_0Output, mb_D_FF700_895MultiplicandStage1Output);

    MB_D_FF_Float_700_895_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF700_895MultiplicandStage1Output, mb_D_FF700_895MultiplicandStage2Output);

    Multiplier_Float_700: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF700_895MultiplicandStage2Output, mb_D_FF700_895MultiplierStage2Output, Multiplier700_Output_895);

    MB_D_FF_Float_Multiplier17_Input2_700_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier697_Output_891, mb_D_FFMultiplier17_Input2_700_0Output);

    MB_D_FF_Float_700_895_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier17_Input2_700_0Output, mb_D_FF700_895MultiplierStage1Output);

    MB_D_FF_Float_700_895_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF700_895MultiplierStage1Output, mb_D_FF700_895MultiplierStage2Output);

    MBRightSHR_Float_701_896: entity work.MBRightSHR(rtl)
    GENERIC MAP (4, NumberOfBits)
    PORT MAP (clk, rst, Multiplier701Weight, mbRightSHR701_896Output);

    MB_D_FF_Float_701_896_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR701_896Output, Multiplier701WeightOutput);

    InputIEEE_Float_701_896: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier701WeightOutput, flopocoMultiplier701WeightOutput);

    MB_D_FF_Float_701_896_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier701WeightOutput, flopocoMultiplier701WeightInput);

    Multiplier_Float_701: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier701WeightInput, mb_D_FF701_896MultiplierStage2Output, Multiplier701_Output_896);

    MB_D_FF_Float_Multiplier21_701_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier21_701_0Input, mb_D_FFMultiplier21_701_0Output);

    MB_D_FF_Float_701_896_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier21_701_0Output, mb_D_FF701_896MultiplierStage1Output);

    MB_D_FF_Float_701_896_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF701_896MultiplierStage1Output, mb_D_FF701_896MultiplierStage2Output);

    MBRightSHR_Float_702_897: entity work.MBRightSHR(rtl)
    GENERIC MAP (4, NumberOfBits)
    PORT MAP (clk, rst, Multiplier702Weight, mbRightSHR702_897Output);

    MB_D_FF_Float_702_897_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR702_897Output, Multiplier702WeightOutput);

    InputIEEE_Float_702_897: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier702WeightOutput, flopocoMultiplier702WeightOutput);

    MB_D_FF_Float_702_897_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier702WeightOutput, flopocoMultiplier702WeightInput);

    Multiplier_Float_702: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier702WeightInput, mb_D_FF702_897MultiplierStage2Output, Multiplier702_Output_897);

    MB_D_FF_Float_Multiplier21_702_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier21_702_0Input, mb_D_FFMultiplier21_702_0Output);

    MB_D_FF_Float_702_897_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier21_702_0Output, mb_D_FF702_897MultiplierStage1Output);

    MB_D_FF_Float_702_897_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF702_897MultiplierStage1Output, mb_D_FF702_897MultiplierStage2Output);

    MB_D_FF_Float_Adder20_Input1_195_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier702_Output_897, mb_D_FFAdder20_Input1_195_0Output);

    MB_D_FF_Float_195_898_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder20_Input1_195_0Output, mb_D_FF195_898AugendStage1Output);

    MB_D_FF_Float_195_898_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF195_898AugendStage1Output, mb_D_FF195_898AugendStage2Output);

    Adder_Float_195: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF195_898AugendStage2Output, mb_D_FF195_898AddendStage2Output, Adder195_Output_898);

    MB_D_FF_Float_Adder20_Input2_195_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier701_Output_896, mb_D_FFAdder20_Input2_195_0Output);

    MB_D_FF_Float_195_898_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder20_Input2_195_0Output, mb_D_FF195_898AddendStage1Output);

    MB_D_FF_Float_195_898_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF195_898AddendStage1Output, mb_D_FF195_898AddendStage2Output);

    MB_D_FF_Float_Multiplier19_703_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder195_Output_898, mb_D_FFMultiplier19_703_0Output);

    MB_D_FF_Float_703_899_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier19_703_0Output, mb_D_FF703_899MultiplierStage1Output);

    MB_D_FF_Float_703_899_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF703_899MultiplierStage1Output, mb_D_FF703_899MultiplierStage2Output);

    Multiplier_Float_703: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF703_899MultiplierStage2Output, mb_D_FF703_899MultiplicandStage2Output, Multiplier703_Output_899);

    MBRightSHR_Float_703_899: entity work.MBRightSHR(rtl)
    GENERIC MAP (36, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR703_899Input, mbRightSHR703_899Output);

    MB_D_FF_Float_703_899_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR703_899Output, mb_D_FF703_899MultiplicandStage1Output);

    MB_D_FF_Float_703_899_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF703_899MultiplicandStage1Output, mb_D_FF703_899MultiplicandStage2Output);

    MB_D_FF_Float_Multiplier18_704_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier703_Output_899, mb_D_FFMultiplier18_704_0Output);

    MB_D_FF_Float_704_900_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier18_704_0Output, mb_D_FF704_900MultiplierStage1Output);

    MB_D_FF_Float_704_900_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF704_900MultiplierStage1Output, mb_D_FF704_900MultiplierStage2Output);

    Multiplier_Float_704: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF704_900MultiplierStage2Output, flopocoMultiplier704WeightInput, Multiplier704_Output_900);

    MBRightSHR_Float_704_900: entity work.MBRightSHR(rtl)
    GENERIC MAP (43, NumberOfBits)
    PORT MAP (clk, rst, Multiplier704Weight, mbRightSHR704_900Output);

    MB_D_FF_Float_704_900_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR704_900Output, Multiplier704WeightOutput);

    InputIEEE_Float_704_900: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier704WeightOutput, flopocoMultiplier704WeightOutput);

    MB_D_FF_Float_704_900_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier704WeightOutput, flopocoMultiplier704WeightInput);

    MB_D_FF_Float_Multiplier17_Input1_707_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder31_Output_165, mb_D_FFMultiplier17_Input1_707_0Output);

    MB_D_FF_Float_707_904_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier17_Input1_707_0Output, mb_D_FF707_904MultiplicandStage1Output);

    MB_D_FF_Float_707_904_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF707_904MultiplicandStage1Output, mb_D_FF707_904MultiplicandStage2Output);

    Multiplier_Float_707: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF707_904MultiplicandStage2Output, mb_D_FF707_904MultiplierStage2Output, Multiplier707_Output_904);

    MB_D_FF_Float_Multiplier17_Input2_707_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier704_Output_900, mb_D_FFMultiplier17_Input2_707_0Output);

    MB_D_FF_Float_707_904_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier17_Input2_707_0Output, mb_D_FF707_904MultiplierStage1Output);

    MB_D_FF_Float_707_904_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF707_904MultiplierStage1Output, mb_D_FF707_904MultiplierStage2Output);

    MB_D_FF_Float_Adder16_Input1_197_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier707_Output_904, mb_D_FFAdder16_Input1_197_0Output);

    MB_D_FF_Float_197_905_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder16_Input1_197_0Output, mb_D_FF197_905AugendStage1Output);

    MB_D_FF_Float_197_905_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF197_905AugendStage1Output, mb_D_FF197_905AugendStage2Output);

    Adder_Float_197: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF197_905AugendStage2Output, mb_D_FF197_905AddendStage2Output, Adder197_Output_905);

    MB_D_FF_Float_Adder16_Input2_197_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier700_Output_895, mb_D_FFAdder16_Input2_197_0Output);

    MB_D_FF_Float_197_905_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder16_Input2_197_0Output, mb_D_FF197_905AddendStage1Output);

    MB_D_FF_Float_197_905_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF197_905AddendStage1Output, mb_D_FF197_905AddendStage2Output);

    MB_D_FF_Float_Multiplier15_708_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder197_Output_905, mb_D_FFMultiplier15_708_0Output);

    MB_D_FF_Float_708_906_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier15_708_0Output, mb_D_FF708_906MultiplierStage1Output);

    MB_D_FF_Float_708_906_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF708_906MultiplierStage1Output, mb_D_FF708_906MultiplierStage2Output);

    Multiplier_Float_708: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF708_906MultiplierStage2Output, mb_D_FF708_906MultiplicandStage2Output, Multiplier708_Output_906);

    MBRightSHR_Float_708_906: entity work.MBRightSHR(rtl)
    GENERIC MAP (82, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR708_906Input, mbRightSHR708_906Output);

    MB_D_FF_Float_708_906_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR708_906Output, mb_D_FF708_906MultiplicandStage1Output);

    MB_D_FF_Float_708_906_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF708_906MultiplicandStage1Output, mb_D_FF708_906MultiplicandStage2Output);

    MB_D_FF_Float_Multiplier14_709_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier708_Output_906, mb_D_FFMultiplier14_709_0Output);

    MB_D_FF_Float_709_907_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier14_709_0Output, mb_D_FF709_907MultiplierStage1Output);

    MB_D_FF_Float_709_907_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF709_907MultiplierStage1Output, mb_D_FF709_907MultiplierStage2Output);

    Multiplier_Float_709: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF709_907MultiplierStage2Output, flopocoMultiplier709WeightInput, Multiplier709_Output_907);

    MBRightSHR_Float_709_907: entity work.MBRightSHR(rtl)
    GENERIC MAP (89, NumberOfBits)
    PORT MAP (clk, rst, Multiplier709Weight, mbRightSHR709_907Output);

    MB_D_FF_Float_709_907_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR709_907Output, Multiplier709WeightOutput);

    InputIEEE_Float_709_907: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier709WeightOutput, flopocoMultiplier709WeightOutput);

    MB_D_FF_Float_709_907_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier709WeightOutput, flopocoMultiplier709WeightInput);

    MB_D_FF_Float_Adder13_Input1_198_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier709_Output_907, mb_D_FFAdder13_Input1_198_0Output);

    MB_D_FF_Float_198_908_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder13_Input1_198_0Output, mb_D_FF198_908AugendStage1Output);

    MB_D_FF_Float_198_908_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF198_908AugendStage1Output, mb_D_FF198_908AugendStage2Output);

    Adder_Float_198: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF198_908AugendStage2Output, mb_D_FF198_908AddendStage2Output, Adder198_Output_908);

    MB_D_FF_Float_Adder13_Input2_198_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier693_Output_886, mb_D_FFAdder13_Input2_198_0Output);

    MB_D_FF_Float_198_908_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder13_Input2_198_0Output, mb_D_FF198_908AddendStage1Output);

    MB_D_FF_Float_198_908_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF198_908AddendStage1Output, mb_D_FF198_908AddendStage2Output);

    MB_D_FF_Float_Multiplier12_710_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder198_Output_908, mb_D_FFMultiplier12_710_0Output);

    MB_D_FF_Float_710_909_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier12_710_0Output, mb_D_FF710_909MultiplierStage1Output);

    MB_D_FF_Float_710_909_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF710_909MultiplierStage1Output, mb_D_FF710_909MultiplierStage2Output);

    Multiplier_Float_710: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF710_909MultiplierStage2Output, mb_D_FF710_909MultiplicandStage2Output, Multiplier710_Output_909);

    MBRightSHR_Float_710_909: entity work.MBRightSHR(rtl)
    GENERIC MAP (121, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR710_909Input, mbRightSHR710_909Output);

    MB_D_FF_Float_710_909_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR710_909Output, mb_D_FF710_909MultiplicandStage1Output);

    MB_D_FF_Float_710_909_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF710_909MultiplicandStage1Output, mb_D_FF710_909MultiplicandStage2Output);

    MB_D_FF_Float_Multiplier11_Input1_721_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder36_Output_184, mb_D_FFMultiplier11_Input1_721_0Output);

    MB_D_FF_Float_721_923_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier11_Input1_721_0Output, mb_D_FF721_923MultiplicandStage1Output);

    MB_D_FF_Float_721_923_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF721_923MultiplicandStage1Output, mb_D_FF721_923MultiplicandStage2Output);

    Multiplier_Float_721: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF721_923MultiplicandStage2Output, mb_D_FF721_923MultiplierStage2Output, Multiplier721_Output_923);

    MB_D_FF_Float_Multiplier11_Input2_721_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier710_Output_909, mb_D_FFMultiplier11_Input2_721_0Output);

    MB_D_FF_Float_721_923_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier11_Input2_721_0Output, mb_D_FF721_923MultiplierStage1Output);

    MB_D_FF_Float_721_923_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF721_923MultiplierStage1Output, mb_D_FF721_923MultiplierStage2Output);

    MB_D_FF_Float_Multiplier14_737_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier692_Output_885, mb_D_FFMultiplier14_737_0Output);

    MB_D_FF_Float_737_944_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier14_737_0Output, mb_D_FF737_944MultiplierStage1Output);

    MB_D_FF_Float_737_944_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF737_944MultiplierStage1Output, mb_D_FF737_944MultiplierStage2Output);

    Multiplier_Float_737: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF737_944MultiplierStage2Output, flopocoMultiplier737WeightInput, Multiplier737_Output_944);

    MBRightSHR_Float_737_944: entity work.MBRightSHR(rtl)
    GENERIC MAP (89, NumberOfBits)
    PORT MAP (clk, rst, Multiplier737Weight, mbRightSHR737_944Output);

    MB_D_FF_Float_737_944_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR737_944Output, Multiplier737WeightOutput);

    InputIEEE_Float_737_944: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier737WeightOutput, flopocoMultiplier737WeightOutput);

    MB_D_FF_Float_737_944_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier737WeightOutput, flopocoMultiplier737WeightInput);

    MB_D_FF_Float_Multiplier14_753_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier708_Output_906, mb_D_FFMultiplier14_753_0Output);

    MB_D_FF_Float_753_965_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier14_753_0Output, mb_D_FF753_965MultiplierStage1Output);

    MB_D_FF_Float_753_965_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF753_965MultiplierStage1Output, mb_D_FF753_965MultiplierStage2Output);

    Multiplier_Float_753: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF753_965MultiplierStage2Output, flopocoMultiplier753WeightInput, Multiplier753_Output_965);

    MBRightSHR_Float_753_965: entity work.MBRightSHR(rtl)
    GENERIC MAP (89, NumberOfBits)
    PORT MAP (clk, rst, Multiplier753Weight, mbRightSHR753_965Output);

    MB_D_FF_Float_753_965_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR753_965Output, Multiplier753WeightOutput);

    InputIEEE_Float_753_965: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier753WeightOutput, flopocoMultiplier753WeightOutput);

    MB_D_FF_Float_753_965_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier753WeightOutput, flopocoMultiplier753WeightInput);

    MB_D_FF_Float_Adder13_Input1_212_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier753_Output_965, mb_D_FFAdder13_Input1_212_0Output);

    MB_D_FF_Float_212_966_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder13_Input1_212_0Output, mb_D_FF212_966AugendStage1Output);

    MB_D_FF_Float_212_966_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF212_966AugendStage1Output, mb_D_FF212_966AugendStage2Output);

    Adder_Float_212: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF212_966AugendStage2Output, mb_D_FF212_966AddendStage2Output, Adder212_Output_966);

    MB_D_FF_Float_Adder13_Input2_212_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier737_Output_944, mb_D_FFAdder13_Input2_212_0Output);

    MB_D_FF_Float_212_966_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder13_Input2_212_0Output, mb_D_FF212_966AddendStage1Output);

    MB_D_FF_Float_212_966_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF212_966AddendStage1Output, mb_D_FF212_966AddendStage2Output);

    MB_D_FF_Float_Multiplier12_754_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder212_Output_966, mb_D_FFMultiplier12_754_0Output);

    MB_D_FF_Float_754_967_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier12_754_0Output, mb_D_FF754_967MultiplierStage1Output);

    MB_D_FF_Float_754_967_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF754_967MultiplierStage1Output, mb_D_FF754_967MultiplierStage2Output);

    Multiplier_Float_754: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF754_967MultiplierStage2Output, mb_D_FF754_967MultiplicandStage2Output, Multiplier754_Output_967);

    MBRightSHR_Float_754_967: entity work.MBRightSHR(rtl)
    GENERIC MAP (121, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR754_967Input, mbRightSHR754_967Output);

    MB_D_FF_Float_754_967_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR754_967Output, mb_D_FF754_967MultiplicandStage1Output);

    MB_D_FF_Float_754_967_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF754_967MultiplicandStage1Output, mb_D_FF754_967MultiplicandStage2Output);

    MB_D_FF_Float_Multiplier11_Input1_765_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder50_Output_242, mb_D_FFMultiplier11_Input1_765_0Output);

    MB_D_FF_Float_765_981_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier11_Input1_765_0Output, mb_D_FF765_981MultiplicandStage1Output);

    MB_D_FF_Float_765_981_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF765_981MultiplicandStage1Output, mb_D_FF765_981MultiplicandStage2Output);

    Multiplier_Float_765: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF765_981MultiplicandStage2Output, mb_D_FF765_981MultiplierStage2Output, Multiplier765_Output_981);

    MB_D_FF_Float_Multiplier11_Input2_765_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier754_Output_967, mb_D_FFMultiplier11_Input2_765_0Output);

    MB_D_FF_Float_765_981_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier11_Input2_765_0Output, mb_D_FF765_981MultiplierStage1Output);

    MB_D_FF_Float_765_981_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF765_981MultiplierStage1Output, mb_D_FF765_981MultiplierStage2Output);

    MB_D_FF_Float_Adder10_Input1_216_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier765_Output_981, mb_D_FFAdder10_Input1_216_0Output);

    MB_D_FF_Float_216_982_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder10_Input1_216_0Output, mb_D_FF216_982AugendStage1Output);

    MB_D_FF_Float_216_982_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF216_982AugendStage1Output, mb_D_FF216_982AugendStage2Output);

    Adder_Float_216: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF216_982AugendStage2Output, mb_D_FF216_982AddendStage2Output, Adder216_Output_982);

    MB_D_FF_Float_Adder10_Input2_216_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier721_Output_923, mb_D_FFAdder10_Input2_216_0Output);

    MB_D_FF_Float_216_982_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder10_Input2_216_0Output, mb_D_FF216_982AddendStage1Output);

    MB_D_FF_Float_216_982_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF216_982AddendStage1Output, mb_D_FF216_982AddendStage2Output);

    MB_D_FF_Float_Multiplier9_766_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder216_Output_982, mb_D_FFMultiplier9_766_0Output);

    MB_D_FF_Float_766_983_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier9_766_0Output, mb_D_FF766_983MultiplierStage1Output);

    MB_D_FF_Float_766_983_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF766_983MultiplierStage1Output, mb_D_FF766_983MultiplierStage2Output);

    Multiplier_Float_766: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF766_983MultiplierStage2Output, mb_D_FF766_983MultiplicandStage2Output, Multiplier766_Output_983);

    MBRightSHR_Float_766_983: entity work.MBRightSHR(rtl)
    GENERIC MAP (160, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR766_983Input, mbRightSHR766_983Output);

    MB_D_FF_Float_766_983_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR766_983Output, mb_D_FF766_983MultiplicandStage1Output);

    MB_D_FF_Float_766_983_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF766_983MultiplicandStage1Output, mb_D_FF766_983MultiplicandStage2Output);

    MB_D_FF_Float_Multiplier8_767_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier766_Output_983, mb_D_FFMultiplier8_767_0Output);

    MB_D_FF_Float_767_984_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier8_767_0Output, mb_D_FF767_984MultiplierStage1Output);

    MB_D_FF_Float_767_984_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF767_984MultiplierStage1Output, mb_D_FF767_984MultiplierStage2Output);

    Multiplier_Float_767: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF767_984MultiplierStage2Output, flopocoMultiplier767WeightInput, Multiplier767_Output_984);

    MBRightSHR_Float_767_984: entity work.MBRightSHR(rtl)
    GENERIC MAP (167, NumberOfBits)
    PORT MAP (clk, rst, Multiplier767Weight, mbRightSHR767_984Output);

    MB_D_FF_Float_767_984_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR767_984Output, Multiplier767WeightOutput);

    InputIEEE_Float_767_984: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier767WeightOutput, flopocoMultiplier767WeightOutput);

    MB_D_FF_Float_767_984_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier767WeightOutput, flopocoMultiplier767WeightInput);

    MB_D_FF_Float_Multiplier17_Input1_774_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder53_Output_254, mb_D_FFMultiplier17_Input1_774_0Output);

    MB_D_FF_Float_774_993_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier17_Input1_774_0Output, mb_D_FF774_993MultiplicandStage1Output);

    MB_D_FF_Float_774_993_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF774_993MultiplicandStage1Output, mb_D_FF774_993MultiplicandStage2Output);

    Multiplier_Float_774: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF774_993MultiplicandStage2Output, mb_D_FF774_993MultiplierStage2Output, Multiplier774_Output_993);

    MB_D_FF_Float_Multiplier17_Input2_774_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier681_Output_870, mb_D_FFMultiplier17_Input2_774_0Output);

    MB_D_FF_Float_774_993_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier17_Input2_774_0Output, mb_D_FF774_993MultiplierStage1Output);

    MB_D_FF_Float_774_993_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF774_993MultiplierStage1Output, mb_D_FF774_993MultiplierStage2Output);

    MB_D_FF_Float_Multiplier17_Input1_781_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder55_Output_263, mb_D_FFMultiplier17_Input1_781_0Output);

    MB_D_FF_Float_781_1002_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier17_Input1_781_0Output, mb_D_FF781_1002MultiplicandStage1Output);

    MB_D_FF_Float_781_1002_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF781_1002MultiplicandStage1Output, mb_D_FF781_1002MultiplicandStage2Output);

    Multiplier_Float_781: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF781_1002MultiplicandStage2Output, mb_D_FF781_1002MultiplierStage2Output, Multiplier781_Output_1002);

    MB_D_FF_Float_Multiplier17_Input2_781_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier688_Output_879, mb_D_FFMultiplier17_Input2_781_0Output);

    MB_D_FF_Float_781_1002_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier17_Input2_781_0Output, mb_D_FF781_1002MultiplierStage1Output);

    MB_D_FF_Float_781_1002_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF781_1002MultiplierStage1Output, mb_D_FF781_1002MultiplierStage2Output);

    MB_D_FF_Float_Adder16_Input1_221_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier781_Output_1002, mb_D_FFAdder16_Input1_221_0Output);

    MB_D_FF_Float_221_1003_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder16_Input1_221_0Output, mb_D_FF221_1003AugendStage1Output);

    MB_D_FF_Float_221_1003_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF221_1003AugendStage1Output, mb_D_FF221_1003AugendStage2Output);

    Adder_Float_221: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF221_1003AugendStage2Output, mb_D_FF221_1003AddendStage2Output, Adder221_Output_1003);

    MB_D_FF_Float_Adder16_Input2_221_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier774_Output_993, mb_D_FFAdder16_Input2_221_0Output);

    MB_D_FF_Float_221_1003_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder16_Input2_221_0Output, mb_D_FF221_1003AddendStage1Output);

    MB_D_FF_Float_221_1003_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF221_1003AddendStage1Output, mb_D_FF221_1003AddendStage2Output);

    MB_D_FF_Float_Multiplier15_782_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder221_Output_1003, mb_D_FFMultiplier15_782_0Output);

    MB_D_FF_Float_782_1004_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier15_782_0Output, mb_D_FF782_1004MultiplierStage1Output);

    MB_D_FF_Float_782_1004_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF782_1004MultiplierStage1Output, mb_D_FF782_1004MultiplierStage2Output);

    Multiplier_Float_782: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF782_1004MultiplierStage2Output, mb_D_FF782_1004MultiplicandStage2Output, Multiplier782_Output_1004);

    MBRightSHR_Float_782_1004: entity work.MBRightSHR(rtl)
    GENERIC MAP (82, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR782_1004Input, mbRightSHR782_1004Output);

    MB_D_FF_Float_782_1004_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR782_1004Output, mb_D_FF782_1004MultiplicandStage1Output);

    MB_D_FF_Float_782_1004_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF782_1004MultiplicandStage1Output, mb_D_FF782_1004MultiplicandStage2Output);

    MB_D_FF_Float_Multiplier14_783_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier782_Output_1004, mb_D_FFMultiplier14_783_0Output);

    MB_D_FF_Float_783_1005_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier14_783_0Output, mb_D_FF783_1005MultiplierStage1Output);

    MB_D_FF_Float_783_1005_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF783_1005MultiplierStage1Output, mb_D_FF783_1005MultiplierStage2Output);

    Multiplier_Float_783: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF783_1005MultiplierStage2Output, flopocoMultiplier783WeightInput, Multiplier783_Output_1005);

    MBRightSHR_Float_783_1005: entity work.MBRightSHR(rtl)
    GENERIC MAP (89, NumberOfBits)
    PORT MAP (clk, rst, Multiplier783Weight, mbRightSHR783_1005Output);

    MB_D_FF_Float_783_1005_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR783_1005Output, Multiplier783WeightOutput);

    InputIEEE_Float_783_1005: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier783WeightOutput, flopocoMultiplier783WeightOutput);

    MB_D_FF_Float_783_1005_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier783WeightOutput, flopocoMultiplier783WeightInput);

    MB_D_FF_Float_Multiplier17_Input1_790_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder58_Output_275, mb_D_FFMultiplier17_Input1_790_0Output);

    MB_D_FF_Float_790_1014_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier17_Input1_790_0Output, mb_D_FF790_1014MultiplicandStage1Output);

    MB_D_FF_Float_790_1014_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF790_1014MultiplicandStage1Output, mb_D_FF790_1014MultiplicandStage2Output);

    Multiplier_Float_790: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF790_1014MultiplicandStage2Output, mb_D_FF790_1014MultiplierStage2Output, Multiplier790_Output_1014);

    MB_D_FF_Float_Multiplier17_Input2_790_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier697_Output_891, mb_D_FFMultiplier17_Input2_790_0Output);

    MB_D_FF_Float_790_1014_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier17_Input2_790_0Output, mb_D_FF790_1014MultiplierStage1Output);

    MB_D_FF_Float_790_1014_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF790_1014MultiplierStage1Output, mb_D_FF790_1014MultiplierStage2Output);

    MB_D_FF_Float_Multiplier17_Input1_797_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder60_Output_284, mb_D_FFMultiplier17_Input1_797_0Output);

    MB_D_FF_Float_797_1023_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier17_Input1_797_0Output, mb_D_FF797_1023MultiplicandStage1Output);

    MB_D_FF_Float_797_1023_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF797_1023MultiplicandStage1Output, mb_D_FF797_1023MultiplicandStage2Output);

    Multiplier_Float_797: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF797_1023MultiplicandStage2Output, mb_D_FF797_1023MultiplierStage2Output, Multiplier797_Output_1023);

    MB_D_FF_Float_Multiplier17_Input2_797_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier704_Output_900, mb_D_FFMultiplier17_Input2_797_0Output);

    MB_D_FF_Float_797_1023_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier17_Input2_797_0Output, mb_D_FF797_1023MultiplierStage1Output);

    MB_D_FF_Float_797_1023_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF797_1023MultiplierStage1Output, mb_D_FF797_1023MultiplierStage2Output);

    MB_D_FF_Float_Adder16_Input1_226_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier797_Output_1023, mb_D_FFAdder16_Input1_226_0Output);

    MB_D_FF_Float_226_1024_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder16_Input1_226_0Output, mb_D_FF226_1024AugendStage1Output);

    MB_D_FF_Float_226_1024_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF226_1024AugendStage1Output, mb_D_FF226_1024AugendStage2Output);

    Adder_Float_226: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF226_1024AugendStage2Output, mb_D_FF226_1024AddendStage2Output, Adder226_Output_1024);

    MB_D_FF_Float_Adder16_Input2_226_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier790_Output_1014, mb_D_FFAdder16_Input2_226_0Output);

    MB_D_FF_Float_226_1024_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder16_Input2_226_0Output, mb_D_FF226_1024AddendStage1Output);

    MB_D_FF_Float_226_1024_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF226_1024AddendStage1Output, mb_D_FF226_1024AddendStage2Output);

    MB_D_FF_Float_Multiplier15_798_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder226_Output_1024, mb_D_FFMultiplier15_798_0Output);

    MB_D_FF_Float_798_1025_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier15_798_0Output, mb_D_FF798_1025MultiplierStage1Output);

    MB_D_FF_Float_798_1025_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF798_1025MultiplierStage1Output, mb_D_FF798_1025MultiplierStage2Output);

    Multiplier_Float_798: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF798_1025MultiplierStage2Output, mb_D_FF798_1025MultiplicandStage2Output, Multiplier798_Output_1025);

    MBRightSHR_Float_798_1025: entity work.MBRightSHR(rtl)
    GENERIC MAP (82, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR798_1025Input, mbRightSHR798_1025Output);

    MB_D_FF_Float_798_1025_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR798_1025Output, mb_D_FF798_1025MultiplicandStage1Output);

    MB_D_FF_Float_798_1025_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF798_1025MultiplicandStage1Output, mb_D_FF798_1025MultiplicandStage2Output);

    MB_D_FF_Float_Multiplier14_799_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier798_Output_1025, mb_D_FFMultiplier14_799_0Output);

    MB_D_FF_Float_799_1026_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier14_799_0Output, mb_D_FF799_1026MultiplierStage1Output);

    MB_D_FF_Float_799_1026_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF799_1026MultiplierStage1Output, mb_D_FF799_1026MultiplierStage2Output);

    Multiplier_Float_799: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF799_1026MultiplierStage2Output, flopocoMultiplier799WeightInput, Multiplier799_Output_1026);

    MBRightSHR_Float_799_1026: entity work.MBRightSHR(rtl)
    GENERIC MAP (89, NumberOfBits)
    PORT MAP (clk, rst, Multiplier799Weight, mbRightSHR799_1026Output);

    MB_D_FF_Float_799_1026_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR799_1026Output, Multiplier799WeightOutput);

    InputIEEE_Float_799_1026: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier799WeightOutput, flopocoMultiplier799WeightOutput);

    MB_D_FF_Float_799_1026_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier799WeightOutput, flopocoMultiplier799WeightInput);

    MB_D_FF_Float_Adder13_Input1_227_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier799_Output_1026, mb_D_FFAdder13_Input1_227_0Output);

    MB_D_FF_Float_227_1027_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder13_Input1_227_0Output, mb_D_FF227_1027AugendStage1Output);

    MB_D_FF_Float_227_1027_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF227_1027AugendStage1Output, mb_D_FF227_1027AugendStage2Output);

    Adder_Float_227: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF227_1027AugendStage2Output, mb_D_FF227_1027AddendStage2Output, Adder227_Output_1027);

    MB_D_FF_Float_Adder13_Input2_227_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier783_Output_1005, mb_D_FFAdder13_Input2_227_0Output);

    MB_D_FF_Float_227_1027_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder13_Input2_227_0Output, mb_D_FF227_1027AddendStage1Output);

    MB_D_FF_Float_227_1027_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF227_1027AddendStage1Output, mb_D_FF227_1027AddendStage2Output);

    MB_D_FF_Float_Multiplier12_800_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder227_Output_1027, mb_D_FFMultiplier12_800_0Output);

    MB_D_FF_Float_800_1028_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier12_800_0Output, mb_D_FF800_1028MultiplierStage1Output);

    MB_D_FF_Float_800_1028_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF800_1028MultiplierStage1Output, mb_D_FF800_1028MultiplierStage2Output);

    Multiplier_Float_800: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF800_1028MultiplierStage2Output, mb_D_FF800_1028MultiplicandStage2Output, Multiplier800_Output_1028);

    MBRightSHR_Float_800_1028: entity work.MBRightSHR(rtl)
    GENERIC MAP (121, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR800_1028Input, mbRightSHR800_1028Output);

    MB_D_FF_Float_800_1028_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR800_1028Output, mb_D_FF800_1028MultiplicandStage1Output);

    MB_D_FF_Float_800_1028_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF800_1028MultiplicandStage1Output, mb_D_FF800_1028MultiplicandStage2Output);

    MB_D_FF_Float_Multiplier11_Input1_811_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder65_Output_303, mb_D_FFMultiplier11_Input1_811_0Output);

    MB_D_FF_Float_811_1042_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier11_Input1_811_0Output, mb_D_FF811_1042MultiplicandStage1Output);

    MB_D_FF_Float_811_1042_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF811_1042MultiplicandStage1Output, mb_D_FF811_1042MultiplicandStage2Output);

    Multiplier_Float_811: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF811_1042MultiplicandStage2Output, mb_D_FF811_1042MultiplierStage2Output, Multiplier811_Output_1042);

    MB_D_FF_Float_Multiplier11_Input2_811_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier800_Output_1028, mb_D_FFMultiplier11_Input2_811_0Output);

    MB_D_FF_Float_811_1042_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier11_Input2_811_0Output, mb_D_FF811_1042MultiplierStage1Output);

    MB_D_FF_Float_811_1042_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF811_1042MultiplierStage1Output, mb_D_FF811_1042MultiplierStage2Output);

    MB_D_FF_Float_Multiplier14_827_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier782_Output_1004, mb_D_FFMultiplier14_827_0Output);

    MB_D_FF_Float_827_1063_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier14_827_0Output, mb_D_FF827_1063MultiplierStage1Output);

    MB_D_FF_Float_827_1063_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF827_1063MultiplierStage1Output, mb_D_FF827_1063MultiplierStage2Output);

    Multiplier_Float_827: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF827_1063MultiplierStage2Output, flopocoMultiplier827WeightInput, Multiplier827_Output_1063);

    MBRightSHR_Float_827_1063: entity work.MBRightSHR(rtl)
    GENERIC MAP (89, NumberOfBits)
    PORT MAP (clk, rst, Multiplier827Weight, mbRightSHR827_1063Output);

    MB_D_FF_Float_827_1063_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR827_1063Output, Multiplier827WeightOutput);

    InputIEEE_Float_827_1063: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier827WeightOutput, flopocoMultiplier827WeightOutput);

    MB_D_FF_Float_827_1063_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier827WeightOutput, flopocoMultiplier827WeightInput);

    MB_D_FF_Float_Multiplier14_843_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier798_Output_1025, mb_D_FFMultiplier14_843_0Output);

    MB_D_FF_Float_843_1084_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier14_843_0Output, mb_D_FF843_1084MultiplierStage1Output);

    MB_D_FF_Float_843_1084_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF843_1084MultiplierStage1Output, mb_D_FF843_1084MultiplierStage2Output);

    Multiplier_Float_843: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF843_1084MultiplierStage2Output, flopocoMultiplier843WeightInput, Multiplier843_Output_1084);

    MBRightSHR_Float_843_1084: entity work.MBRightSHR(rtl)
    GENERIC MAP (89, NumberOfBits)
    PORT MAP (clk, rst, Multiplier843Weight, mbRightSHR843_1084Output);

    MB_D_FF_Float_843_1084_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR843_1084Output, Multiplier843WeightOutput);

    InputIEEE_Float_843_1084: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier843WeightOutput, flopocoMultiplier843WeightOutput);

    MB_D_FF_Float_843_1084_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier843WeightOutput, flopocoMultiplier843WeightInput);

    MB_D_FF_Float_Adder13_Input1_241_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier843_Output_1084, mb_D_FFAdder13_Input1_241_0Output);

    MB_D_FF_Float_241_1085_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder13_Input1_241_0Output, mb_D_FF241_1085AugendStage1Output);

    MB_D_FF_Float_241_1085_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF241_1085AugendStage1Output, mb_D_FF241_1085AugendStage2Output);

    Adder_Float_241: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF241_1085AugendStage2Output, mb_D_FF241_1085AddendStage2Output, Adder241_Output_1085);

    MB_D_FF_Float_Adder13_Input2_241_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier827_Output_1063, mb_D_FFAdder13_Input2_241_0Output);

    MB_D_FF_Float_241_1085_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder13_Input2_241_0Output, mb_D_FF241_1085AddendStage1Output);

    MB_D_FF_Float_241_1085_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF241_1085AddendStage1Output, mb_D_FF241_1085AddendStage2Output);

    MB_D_FF_Float_Multiplier12_844_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder241_Output_1085, mb_D_FFMultiplier12_844_0Output);

    MB_D_FF_Float_844_1086_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier12_844_0Output, mb_D_FF844_1086MultiplierStage1Output);

    MB_D_FF_Float_844_1086_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF844_1086MultiplierStage1Output, mb_D_FF844_1086MultiplierStage2Output);

    Multiplier_Float_844: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF844_1086MultiplierStage2Output, mb_D_FF844_1086MultiplicandStage2Output, Multiplier844_Output_1086);

    MBRightSHR_Float_844_1086: entity work.MBRightSHR(rtl)
    GENERIC MAP (121, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR844_1086Input, mbRightSHR844_1086Output);

    MB_D_FF_Float_844_1086_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR844_1086Output, mb_D_FF844_1086MultiplicandStage1Output);

    MB_D_FF_Float_844_1086_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF844_1086MultiplicandStage1Output, mb_D_FF844_1086MultiplicandStage2Output);

    MB_D_FF_Float_Multiplier11_Input1_855_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder79_Output_361, mb_D_FFMultiplier11_Input1_855_0Output);

    MB_D_FF_Float_855_1100_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier11_Input1_855_0Output, mb_D_FF855_1100MultiplicandStage1Output);

    MB_D_FF_Float_855_1100_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF855_1100MultiplicandStage1Output, mb_D_FF855_1100MultiplicandStage2Output);

    Multiplier_Float_855: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF855_1100MultiplicandStage2Output, mb_D_FF855_1100MultiplierStage2Output, Multiplier855_Output_1100);

    MB_D_FF_Float_Multiplier11_Input2_855_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier844_Output_1086, mb_D_FFMultiplier11_Input2_855_0Output);

    MB_D_FF_Float_855_1100_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier11_Input2_855_0Output, mb_D_FF855_1100MultiplierStage1Output);

    MB_D_FF_Float_855_1100_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF855_1100MultiplierStage1Output, mb_D_FF855_1100MultiplierStage2Output);

    MB_D_FF_Float_Adder10_Input1_245_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier855_Output_1100, mb_D_FFAdder10_Input1_245_0Output);

    MB_D_FF_Float_245_1101_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder10_Input1_245_0Output, mb_D_FF245_1101AugendStage1Output);

    MB_D_FF_Float_245_1101_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF245_1101AugendStage1Output, mb_D_FF245_1101AugendStage2Output);

    Adder_Float_245: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF245_1101AugendStage2Output, mb_D_FF245_1101AddendStage2Output, Adder245_Output_1101);

    MB_D_FF_Float_Adder10_Input2_245_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier811_Output_1042, mb_D_FFAdder10_Input2_245_0Output);

    MB_D_FF_Float_245_1101_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder10_Input2_245_0Output, mb_D_FF245_1101AddendStage1Output);

    MB_D_FF_Float_245_1101_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF245_1101AddendStage1Output, mb_D_FF245_1101AddendStage2Output);

    MB_D_FF_Float_Multiplier9_856_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder245_Output_1101, mb_D_FFMultiplier9_856_0Output);

    MB_D_FF_Float_856_1102_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier9_856_0Output, mb_D_FF856_1102MultiplierStage1Output);

    MB_D_FF_Float_856_1102_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF856_1102MultiplierStage1Output, mb_D_FF856_1102MultiplierStage2Output);

    Multiplier_Float_856: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF856_1102MultiplierStage2Output, mb_D_FF856_1102MultiplicandStage2Output, Multiplier856_Output_1102);

    MBRightSHR_Float_856_1102: entity work.MBRightSHR(rtl)
    GENERIC MAP (160, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR856_1102Input, mbRightSHR856_1102Output);

    MB_D_FF_Float_856_1102_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR856_1102Output, mb_D_FF856_1102MultiplicandStage1Output);

    MB_D_FF_Float_856_1102_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF856_1102MultiplicandStage1Output, mb_D_FF856_1102MultiplicandStage2Output);

    MB_D_FF_Float_Multiplier8_857_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier856_Output_1102, mb_D_FFMultiplier8_857_0Output);

    MB_D_FF_Float_857_1103_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier8_857_0Output, mb_D_FF857_1103MultiplierStage1Output);

    MB_D_FF_Float_857_1103_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF857_1103MultiplierStage1Output, mb_D_FF857_1103MultiplierStage2Output);

    Multiplier_Float_857: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF857_1103MultiplierStage2Output, flopocoMultiplier857WeightInput, Multiplier857_Output_1103);

    MBRightSHR_Float_857_1103: entity work.MBRightSHR(rtl)
    GENERIC MAP (167, NumberOfBits)
    PORT MAP (clk, rst, Multiplier857Weight, mbRightSHR857_1103Output);

    MB_D_FF_Float_857_1103_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR857_1103Output, Multiplier857WeightOutput);

    InputIEEE_Float_857_1103: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier857WeightOutput, flopocoMultiplier857WeightOutput);

    MB_D_FF_Float_857_1103_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier857WeightOutput, flopocoMultiplier857WeightInput);

    MB_D_FF_Float_Adder7_Input1_246_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier857_Output_1103, mb_D_FFAdder7_Input1_246_0Output);

    MB_D_FF_Float_246_1104_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder7_Input1_246_0Output, mb_D_FF246_1104AugendStage1Output);

    MB_D_FF_Float_246_1104_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF246_1104AugendStage1Output, mb_D_FF246_1104AugendStage2Output);

    Adder_Float_246: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF246_1104AugendStage2Output, mb_D_FF246_1104AddendStage2Output, Adder246_Output_1104);

    MB_D_FF_Float_Adder7_Input2_246_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier767_Output_984, mb_D_FFAdder7_Input2_246_0Output);

    MB_D_FF_Float_246_1104_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder7_Input2_246_0Output, mb_D_FF246_1104AddendStage1Output);

    MB_D_FF_Float_246_1104_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF246_1104AddendStage1Output, mb_D_FF246_1104AddendStage2Output);

    MB_D_FF_Float_Multiplier6_Input1_858_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder246_Output_1104, mb_D_FFMultiplier6_Input1_858_0Output);

    MB_D_FF_Float_858_1105_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier6_Input1_858_0Output, mb_D_FF858_1105MultiplicandStage1Output);

    MB_D_FF_Float_858_1105_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF858_1105MultiplicandStage1Output, mb_D_FF858_1105MultiplicandStage2Output);

    Multiplier_Float_858: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF858_1105MultiplicandStage2Output, mb_D_FF858_1105MultiplierStage2Output, Multiplier858_Output_1105);

    MB_D_FF_Float_Multiplier6_Input2_858_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier677_Output_865, mb_D_FFMultiplier6_Input2_858_0Output);

    MB_D_FF_Float_858_1105_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier6_Input2_858_0Output, mb_D_FF858_1105MultiplierStage1Output);

    MB_D_FF_Float_858_1105_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF858_1105MultiplierStage1Output, mb_D_FF858_1105MultiplierStage2Output);

    MB_D_FF_Float_Multiplier12_883_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier596_Output_766, mb_D_FFMultiplier12_883_0Output);

    MB_D_FF_Float_883_1135_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier12_883_0Output, mb_D_FF883_1135MultiplierStage1Output);

    MB_D_FF_Float_883_1135_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF883_1135MultiplierStage1Output, mb_D_FF883_1135MultiplierStage2Output);

    Multiplier_Float_883: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF883_1135MultiplierStage2Output, flopocoMultiplier883WeightInput, Multiplier883_Output_1135);

    MBRightSHR_Float_883_1135: entity work.MBRightSHR(rtl)
    GENERIC MAP (121, NumberOfBits)
    PORT MAP (clk, rst, Multiplier883Weight, mbRightSHR883_1135Output);

    MB_D_FF_Float_883_1135_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR883_1135Output, Multiplier883WeightOutput);

    InputIEEE_Float_883_1135: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier883WeightOutput, flopocoMultiplier883WeightOutput);

    MB_D_FF_Float_883_1135_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier883WeightOutput, flopocoMultiplier883WeightInput);

    MB_D_FF_Float_Multiplier12_908_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier621_Output_796, mb_D_FFMultiplier12_908_0Output);

    MB_D_FF_Float_908_1165_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier12_908_0Output, mb_D_FF908_1165MultiplierStage1Output);

    MB_D_FF_Float_908_1165_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF908_1165MultiplierStage1Output, mb_D_FF908_1165MultiplierStage2Output);

    Multiplier_Float_908: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF908_1165MultiplierStage2Output, flopocoMultiplier908WeightInput, Multiplier908_Output_1165);

    MBRightSHR_Float_908_1165: entity work.MBRightSHR(rtl)
    GENERIC MAP (121, NumberOfBits)
    PORT MAP (clk, rst, Multiplier908Weight, mbRightSHR908_1165Output);

    MB_D_FF_Float_908_1165_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR908_1165Output, Multiplier908WeightOutput);

    InputIEEE_Float_908_1165: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier908WeightOutput, flopocoMultiplier908WeightOutput);

    MB_D_FF_Float_908_1165_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier908WeightOutput, flopocoMultiplier908WeightInput);

    MB_D_FF_Float_Adder11_Input1_257_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier908_Output_1165, mb_D_FFAdder11_Input1_257_0Output);

    MB_D_FF_Float_257_1166_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder11_Input1_257_0Output, mb_D_FF257_1166AugendStage1Output);

    MB_D_FF_Float_257_1166_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF257_1166AugendStage1Output, mb_D_FF257_1166AugendStage2Output);

    Adder_Float_257: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF257_1166AugendStage2Output, mb_D_FF257_1166AddendStage2Output, Adder257_Output_1166);

    MB_D_FF_Float_Adder11_Input2_257_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier883_Output_1135, mb_D_FFAdder11_Input2_257_0Output);

    MB_D_FF_Float_257_1166_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder11_Input2_257_0Output, mb_D_FF257_1166AddendStage1Output);

    MB_D_FF_Float_257_1166_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF257_1166AddendStage1Output, mb_D_FF257_1166AddendStage2Output);

    MB_D_FF_Float_Multiplier10_909_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder257_Output_1166, mb_D_FFMultiplier10_909_0Output);

    MB_D_FF_Float_909_1167_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier10_909_0Output, mb_D_FF909_1167MultiplierStage1Output);

    MB_D_FF_Float_909_1167_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF909_1167MultiplierStage1Output, mb_D_FF909_1167MultiplierStage2Output);

    Multiplier_Float_909: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF909_1167MultiplierStage2Output, mb_D_FF909_1167MultiplicandStage2Output, Multiplier909_Output_1167);

    MBRightSHR_Float_909_1167: entity work.MBRightSHR(rtl)
    GENERIC MAP (135, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR909_1167Input, mbRightSHR909_1167Output);

    MB_D_FF_Float_909_1167_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR909_1167Output, mb_D_FF909_1167MultiplicandStage1Output);

    MB_D_FF_Float_909_1167_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF909_1167MultiplicandStage1Output, mb_D_FF909_1167MultiplicandStage2Output);

    MB_D_FF_Float_Multiplier9_910_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier909_Output_1167, mb_D_FFMultiplier9_910_0Output);

    MB_D_FF_Float_910_1168_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier9_910_0Output, mb_D_FF910_1168MultiplierStage1Output);

    MB_D_FF_Float_910_1168_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF910_1168MultiplierStage1Output, mb_D_FF910_1168MultiplierStage2Output);

    Multiplier_Float_910: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF910_1168MultiplierStage2Output, flopocoMultiplier910WeightInput, Multiplier910_Output_1168);

    MBRightSHR_Float_910_1168: entity work.MBRightSHR(rtl)
    GENERIC MAP (160, NumberOfBits)
    PORT MAP (clk, rst, Multiplier910Weight, mbRightSHR910_1168Output);

    MB_D_FF_Float_910_1168_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR910_1168Output, Multiplier910WeightOutput);

    InputIEEE_Float_910_1168: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier910WeightOutput, flopocoMultiplier910WeightOutput);

    MB_D_FF_Float_910_1168_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier910WeightOutput, flopocoMultiplier910WeightInput);

    MB_D_FF_Float_Multiplier12_935_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier648_Output_829, mb_D_FFMultiplier12_935_0Output);

    MB_D_FF_Float_935_1198_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier12_935_0Output, mb_D_FF935_1198MultiplierStage1Output);

    MB_D_FF_Float_935_1198_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF935_1198MultiplierStage1Output, mb_D_FF935_1198MultiplierStage2Output);

    Multiplier_Float_935: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF935_1198MultiplierStage2Output, flopocoMultiplier935WeightInput, Multiplier935_Output_1198);

    MBRightSHR_Float_935_1198: entity work.MBRightSHR(rtl)
    GENERIC MAP (121, NumberOfBits)
    PORT MAP (clk, rst, Multiplier935Weight, mbRightSHR935_1198Output);

    MB_D_FF_Float_935_1198_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR935_1198Output, Multiplier935WeightOutput);

    InputIEEE_Float_935_1198: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier935WeightOutput, flopocoMultiplier935WeightOutput);

    MB_D_FF_Float_935_1198_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier935WeightOutput, flopocoMultiplier935WeightInput);

    MB_D_FF_Float_Multiplier12_960_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier673_Output_859, mb_D_FFMultiplier12_960_0Output);

    MB_D_FF_Float_960_1228_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier12_960_0Output, mb_D_FF960_1228MultiplierStage1Output);

    MB_D_FF_Float_960_1228_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF960_1228MultiplierStage1Output, mb_D_FF960_1228MultiplierStage2Output);

    Multiplier_Float_960: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF960_1228MultiplierStage2Output, flopocoMultiplier960WeightInput, Multiplier960_Output_1228);

    MBRightSHR_Float_960_1228: entity work.MBRightSHR(rtl)
    GENERIC MAP (121, NumberOfBits)
    PORT MAP (clk, rst, Multiplier960Weight, mbRightSHR960_1228Output);

    MB_D_FF_Float_960_1228_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR960_1228Output, Multiplier960WeightOutput);

    InputIEEE_Float_960_1228: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier960WeightOutput, flopocoMultiplier960WeightOutput);

    MB_D_FF_Float_960_1228_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier960WeightOutput, flopocoMultiplier960WeightInput);

    MB_D_FF_Float_Adder11_Input1_268_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier960_Output_1228, mb_D_FFAdder11_Input1_268_0Output);

    MB_D_FF_Float_268_1229_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder11_Input1_268_0Output, mb_D_FF268_1229AugendStage1Output);

    MB_D_FF_Float_268_1229_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF268_1229AugendStage1Output, mb_D_FF268_1229AugendStage2Output);

    Adder_Float_268: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF268_1229AugendStage2Output, mb_D_FF268_1229AddendStage2Output, Adder268_Output_1229);

    MB_D_FF_Float_Adder11_Input2_268_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier935_Output_1198, mb_D_FFAdder11_Input2_268_0Output);

    MB_D_FF_Float_268_1229_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder11_Input2_268_0Output, mb_D_FF268_1229AddendStage1Output);

    MB_D_FF_Float_268_1229_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF268_1229AddendStage1Output, mb_D_FF268_1229AddendStage2Output);

    MB_D_FF_Float_Multiplier10_961_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder268_Output_1229, mb_D_FFMultiplier10_961_0Output);

    MB_D_FF_Float_961_1230_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier10_961_0Output, mb_D_FF961_1230MultiplierStage1Output);

    MB_D_FF_Float_961_1230_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF961_1230MultiplierStage1Output, mb_D_FF961_1230MultiplierStage2Output);

    Multiplier_Float_961: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF961_1230MultiplierStage2Output, mb_D_FF961_1230MultiplicandStage2Output, Multiplier961_Output_1230);

    MBRightSHR_Float_961_1230: entity work.MBRightSHR(rtl)
    GENERIC MAP (135, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR961_1230Input, mbRightSHR961_1230Output);

    MB_D_FF_Float_961_1230_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR961_1230Output, mb_D_FF961_1230MultiplicandStage1Output);

    MB_D_FF_Float_961_1230_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF961_1230MultiplicandStage1Output, mb_D_FF961_1230MultiplicandStage2Output);

    MB_D_FF_Float_Multiplier9_962_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier961_Output_1230, mb_D_FFMultiplier9_962_0Output);

    MB_D_FF_Float_962_1231_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier9_962_0Output, mb_D_FF962_1231MultiplierStage1Output);

    MB_D_FF_Float_962_1231_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF962_1231MultiplierStage1Output, mb_D_FF962_1231MultiplierStage2Output);

    Multiplier_Float_962: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF962_1231MultiplierStage2Output, flopocoMultiplier962WeightInput, Multiplier962_Output_1231);

    MBRightSHR_Float_962_1231: entity work.MBRightSHR(rtl)
    GENERIC MAP (160, NumberOfBits)
    PORT MAP (clk, rst, Multiplier962Weight, mbRightSHR962_1231Output);

    MB_D_FF_Float_962_1231_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR962_1231Output, Multiplier962WeightOutput);

    InputIEEE_Float_962_1231: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier962WeightOutput, flopocoMultiplier962WeightOutput);

    MB_D_FF_Float_962_1231_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier962WeightOutput, flopocoMultiplier962WeightInput);

    MB_D_FF_Float_Adder8_Input1_269_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier962_Output_1231, mb_D_FFAdder8_Input1_269_0Output);

    MB_D_FF_Float_269_1232_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder8_Input1_269_0Output, mb_D_FF269_1232AugendStage1Output);

    MB_D_FF_Float_269_1232_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF269_1232AugendStage1Output, mb_D_FF269_1232AugendStage2Output);

    Adder_Float_269: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF269_1232AugendStage2Output, mb_D_FF269_1232AddendStage2Output, Adder269_Output_1232);

    MB_D_FF_Float_Adder8_Input2_269_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier910_Output_1168, mb_D_FFAdder8_Input2_269_0Output);

    MB_D_FF_Float_269_1232_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder8_Input2_269_0Output, mb_D_FF269_1232AddendStage1Output);

    MB_D_FF_Float_269_1232_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF269_1232AddendStage1Output, mb_D_FF269_1232AddendStage2Output);

    MB_D_FF_Float_Multiplier7_963_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder269_Output_1232, mb_D_FFMultiplier7_963_0Output);

    MB_D_FF_Float_963_1233_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier7_963_0Output, mb_D_FF963_1233MultiplierStage1Output);

    MB_D_FF_Float_963_1233_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF963_1233MultiplierStage1Output, mb_D_FF963_1233MultiplierStage2Output);

    Multiplier_Float_963: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF963_1233MultiplierStage2Output, mb_D_FF963_1233MultiplicandStage2Output, Multiplier963_Output_1233);

    MBRightSHR_Float_963_1233: entity work.MBRightSHR(rtl)
    GENERIC MAP (174, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR963_1233Input, mbRightSHR963_1233Output);

    MB_D_FF_Float_963_1233_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR963_1233Output, mb_D_FF963_1233MultiplicandStage1Output);

    MB_D_FF_Float_963_1233_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF963_1233MultiplicandStage1Output, mb_D_FF963_1233MultiplicandStage2Output);

    MB_D_FF_Float_Multiplier8_1053_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier766_Output_983, mb_D_FFMultiplier8_1053_0Output);

    MB_D_FF_Float_1053_1352_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier8_1053_0Output, mb_D_FF1053_1352MultiplierStage1Output);

    MB_D_FF_Float_1053_1352_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1053_1352MultiplierStage1Output, mb_D_FF1053_1352MultiplierStage2Output);

    Multiplier_Float_1053: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF1053_1352MultiplierStage2Output, flopocoMultiplier1053WeightInput, Multiplier1053_Output_1352);

    MBRightSHR_Float_1053_1352: entity work.MBRightSHR(rtl)
    GENERIC MAP (167, NumberOfBits)
    PORT MAP (clk, rst, Multiplier1053Weight, mbRightSHR1053_1352Output);

    MB_D_FF_Float_1053_1352_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR1053_1352Output, Multiplier1053WeightOutput);

    InputIEEE_Float_1053_1352: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier1053WeightOutput, flopocoMultiplier1053WeightOutput);

    MB_D_FF_Float_1053_1352_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier1053WeightOutput, flopocoMultiplier1053WeightInput);

    MB_D_FF_Float_Multiplier8_1143_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier856_Output_1102, mb_D_FFMultiplier8_1143_0Output);

    MB_D_FF_Float_1143_1471_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier8_1143_0Output, mb_D_FF1143_1471MultiplierStage1Output);

    MB_D_FF_Float_1143_1471_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1143_1471MultiplierStage1Output, mb_D_FF1143_1471MultiplierStage2Output);

    Multiplier_Float_1143: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF1143_1471MultiplierStage2Output, flopocoMultiplier1143WeightInput, Multiplier1143_Output_1471);

    MBRightSHR_Float_1143_1471: entity work.MBRightSHR(rtl)
    GENERIC MAP (167, NumberOfBits)
    PORT MAP (clk, rst, Multiplier1143Weight, mbRightSHR1143_1471Output);

    MB_D_FF_Float_1143_1471_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR1143_1471Output, Multiplier1143WeightOutput);

    InputIEEE_Float_1143_1471: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier1143WeightOutput, flopocoMultiplier1143WeightOutput);

    MB_D_FF_Float_1143_1471_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier1143WeightOutput, flopocoMultiplier1143WeightInput);

    MB_D_FF_Float_Adder7_Input1_328_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier1143_Output_1471, mb_D_FFAdder7_Input1_328_0Output);

    MB_D_FF_Float_328_1472_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder7_Input1_328_0Output, mb_D_FF328_1472AugendStage1Output);

    MB_D_FF_Float_328_1472_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF328_1472AugendStage1Output, mb_D_FF328_1472AugendStage2Output);

    Adder_Float_328: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF328_1472AugendStage2Output, mb_D_FF328_1472AddendStage2Output, Adder328_Output_1472);

    MB_D_FF_Float_Adder7_Input2_328_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier1053_Output_1352, mb_D_FFAdder7_Input2_328_0Output);

    MB_D_FF_Float_328_1472_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder7_Input2_328_0Output, mb_D_FF328_1472AddendStage1Output);

    MB_D_FF_Float_328_1472_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF328_1472AddendStage1Output, mb_D_FF328_1472AddendStage2Output);

    MB_D_FF_Float_Multiplier6_Input1_1144_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder328_Output_1472, mb_D_FFMultiplier6_Input1_1144_0Output);

    MB_D_FF_Float_1144_1473_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier6_Input1_1144_0Output, mb_D_FF1144_1473MultiplicandStage1Output);

    MB_D_FF_Float_1144_1473_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1144_1473MultiplicandStage1Output, mb_D_FF1144_1473MultiplicandStage2Output);

    Multiplier_Float_1144: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF1144_1473MultiplicandStage2Output, mb_D_FF1144_1473MultiplierStage2Output, Multiplier1144_Output_1473);

    MB_D_FF_Float_Multiplier6_Input2_1144_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier963_Output_1233, mb_D_FFMultiplier6_Input2_1144_0Output);

    MB_D_FF_Float_1144_1473_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier6_Input2_1144_0Output, mb_D_FF1144_1473MultiplierStage1Output);

    MB_D_FF_Float_1144_1473_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1144_1473MultiplierStage1Output, mb_D_FF1144_1473MultiplierStage2Output);

    MB_D_FF_Float_Adder5_Input1_329_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier1144_Output_1473, mb_D_FFAdder5_Input1_329_0Output);

    MB_D_FF_Float_329_1474_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder5_Input1_329_0Output, mb_D_FF329_1474AugendStage1Output);

    MB_D_FF_Float_329_1474_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF329_1474AugendStage1Output, mb_D_FF329_1474AugendStage2Output);

    Adder_Float_329: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF329_1474AugendStage2Output, mb_D_FF329_1474AddendStage2Output, Adder329_Output_1474);

    MB_D_FF_Float_Adder5_Input2_329_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier858_Output_1105, mb_D_FFAdder5_Input2_329_0Output);

    MB_D_FF_Float_329_1474_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder5_Input2_329_0Output, mb_D_FF329_1474AddendStage1Output);

    MB_D_FF_Float_329_1474_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF329_1474AddendStage1Output, mb_D_FF329_1474AddendStage2Output);

    MB_D_FF_Float_Multiplier4_1145_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder329_Output_1474, mb_D_FFMultiplier4_1145_0Output);

    MB_D_FF_Float_1145_1475_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier4_1145_0Output, mb_D_FF1145_1475MultiplierStage1Output);

    MB_D_FF_Float_1145_1475_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1145_1475MultiplierStage1Output, mb_D_FF1145_1475MultiplierStage2Output);

    Multiplier_Float_1145: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF1145_1475MultiplierStage2Output, mb_D_FF1145_1475MultiplicandStage2Output, Multiplier1145_Output_1475);

    MBRightSHR_Float_1145_1475: entity work.MBRightSHR(rtl)
    GENERIC MAP (231, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR1145_1475Input, mbRightSHR1145_1475Output);

    MB_D_FF_Float_1145_1475_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR1145_1475Output, mb_D_FF1145_1475MultiplicandStage1Output);

    MB_D_FF_Float_1145_1475_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1145_1475MultiplicandStage1Output, mb_D_FF1145_1475MultiplicandStage2Output);

    MB_D_FF_Float_Adder3_Input1_330_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier1145_Output_1475, mb_D_FFAdder3_Input1_330_0Output);

    MB_D_FF_Float_330_1476_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder3_Input1_330_0Output, mb_D_FF330_1476AugendStage1Output);

    MB_D_FF_Float_330_1476_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF330_1476AugendStage1Output, mb_D_FF330_1476AugendStage2Output);

    Adder_Float_330: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF330_1476AugendStage2Output, mb_D_FF330_1476AddendStage2Output, Adder330_Output_1476);

    MB_D_FF_Float_Adder3_Input2_330_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier572_Output_737, mb_D_FFAdder3_Input2_330_0Output);

    MB_D_FF_Float_330_1476_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder3_Input2_330_0Output, mb_D_FF330_1476AddendStage1Output);

    MB_D_FF_Float_330_1476_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF330_1476AddendStage1Output, mb_D_FF330_1476AddendStage2Output);

    MB_D_FF_Float_Multiplier2_1146_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder330_Output_1476, mb_D_FFMultiplier2_1146_0Output);

    MB_D_FF_Float_1146_1477_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier2_1146_0Output, mb_D_FF1146_1477MultiplierStage1Output);

    MB_D_FF_Float_1146_1477_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1146_1477MultiplierStage1Output, mb_D_FF1146_1477MultiplierStage2Output);

    Multiplier_Float_1146: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF1146_1477MultiplierStage2Output, mb_D_FF1146_1477MultiplicandStage2Output, Multiplier1146_Output_1477);

    MBRightSHR_Float_1146_1477: entity work.MBRightSHR(rtl)
    GENERIC MAP (263, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR1146_1477Input, mbRightSHR1146_1477Output);

    MB_D_FF_Float_1146_1477_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR1146_1477Output, mb_D_FF1146_1477MultiplicandStage1Output);

    MB_D_FF_Float_1146_1477_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1146_1477MultiplicandStage1Output, mb_D_FF1146_1477MultiplicandStage2Output);

    MB_D_FF_Float_Multiplier9_1198_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier50_Output_61, mb_D_FFMultiplier9_1198_0Output);

    MB_D_FF_Float_1198_1540_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier9_1198_0Output, mb_D_FF1198_1540MultiplierStage1Output);

    MB_D_FF_Float_1198_1540_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1198_1540MultiplierStage1Output, mb_D_FF1198_1540MultiplierStage2Output);

    Multiplier_Float_1198: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF1198_1540MultiplierStage2Output, flopocoMultiplier1198WeightInput, Multiplier1198_Output_1540);

    MBRightSHR_Float_1198_1540: entity work.MBRightSHR(rtl)
    GENERIC MAP (160, NumberOfBits)
    PORT MAP (clk, rst, Multiplier1198Weight, mbRightSHR1198_1540Output);

    MB_D_FF_Float_1198_1540_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR1198_1540Output, Multiplier1198WeightOutput);

    InputIEEE_Float_1198_1540: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier1198WeightOutput, flopocoMultiplier1198WeightOutput);

    MB_D_FF_Float_1198_1540_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier1198WeightOutput, flopocoMultiplier1198WeightInput);

    MB_D_FF_Float_Multiplier9_1250_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier102_Output_124, mb_D_FFMultiplier9_1250_0Output);

    MB_D_FF_Float_1250_1603_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier9_1250_0Output, mb_D_FF1250_1603MultiplierStage1Output);

    MB_D_FF_Float_1250_1603_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1250_1603MultiplierStage1Output, mb_D_FF1250_1603MultiplierStage2Output);

    Multiplier_Float_1250: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF1250_1603MultiplierStage2Output, flopocoMultiplier1250WeightInput, Multiplier1250_Output_1603);

    MBRightSHR_Float_1250_1603: entity work.MBRightSHR(rtl)
    GENERIC MAP (160, NumberOfBits)
    PORT MAP (clk, rst, Multiplier1250Weight, mbRightSHR1250_1603Output);

    MB_D_FF_Float_1250_1603_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR1250_1603Output, Multiplier1250WeightOutput);

    InputIEEE_Float_1250_1603: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier1250WeightOutput, flopocoMultiplier1250WeightOutput);

    MB_D_FF_Float_1250_1603_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier1250WeightOutput, flopocoMultiplier1250WeightInput);

    MB_D_FF_Float_Adder8_Input1_353_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier1250_Output_1603, mb_D_FFAdder8_Input1_353_0Output);

    MB_D_FF_Float_353_1604_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder8_Input1_353_0Output, mb_D_FF353_1604AugendStage1Output);

    MB_D_FF_Float_353_1604_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF353_1604AugendStage1Output, mb_D_FF353_1604AugendStage2Output);

    Adder_Float_353: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF353_1604AugendStage2Output, mb_D_FF353_1604AddendStage2Output, Adder353_Output_1604);

    MB_D_FF_Float_Adder8_Input2_353_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier1198_Output_1540, mb_D_FFAdder8_Input2_353_0Output);

    MB_D_FF_Float_353_1604_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder8_Input2_353_0Output, mb_D_FF353_1604AddendStage1Output);

    MB_D_FF_Float_353_1604_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF353_1604AddendStage1Output, mb_D_FF353_1604AddendStage2Output);

    MB_D_FF_Float_Multiplier7_1251_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder353_Output_1604, mb_D_FFMultiplier7_1251_0Output);

    MB_D_FF_Float_1251_1605_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier7_1251_0Output, mb_D_FF1251_1605MultiplierStage1Output);

    MB_D_FF_Float_1251_1605_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1251_1605MultiplierStage1Output, mb_D_FF1251_1605MultiplierStage2Output);

    Multiplier_Float_1251: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF1251_1605MultiplierStage2Output, mb_D_FF1251_1605MultiplicandStage2Output, Multiplier1251_Output_1605);

    MBRightSHR_Float_1251_1605: entity work.MBRightSHR(rtl)
    GENERIC MAP (174, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR1251_1605Input, mbRightSHR1251_1605Output);

    MB_D_FF_Float_1251_1605_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR1251_1605Output, mb_D_FF1251_1605MultiplicandStage1Output);

    MB_D_FF_Float_1251_1605_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1251_1605MultiplicandStage1Output, mb_D_FF1251_1605MultiplicandStage2Output);

    MBRightSHR_Float_1285_Input11650: entity work.MBRightSHR(rtl)
    GENERIC MAP (50, NumberOfBits)
    PORT MAP (clk, rst, Multiplier1285Weight, mbRightSHR1285_Input1_1650Output);

    MB_D_FF_Float_1285_1650_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR1285_Input1_1650Output, Multiplier1285WeightOutput);

    InputIEEE_Float_1285_1650: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier1285WeightOutput, flopocoMultiplier1285WeightOutput);

    MB_D_FF_Float_1285_1650_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier1285WeightOutput, flopocoMultiplier1285WeightInput);

    Multiplier_Float_1285: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier1285WeightInput, mb_D_FF1285_1650MultiplierStage2Output, Multiplier1285_Output_1650);

    MBRightSHR_Float_1285_Input2_1650: entity work.MBRightSHR(rtl)
    GENERIC MAP (50, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR1285_Input2_1650Input, mbRightSHR1285_Input2_1650Output);

    MB_D_FF_Float_1285_1650_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR1285_Input2_1650Output, mb_D_FF1285_1650MultiplierStage1Output);

    MB_D_FF_Float_1285_1650_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1285_1650MultiplierStage1Output, mb_D_FF1285_1650MultiplierStage2Output);

    MBRightSHR_Float_1286_Input11651: entity work.MBRightSHR(rtl)
    GENERIC MAP (50, NumberOfBits)
    PORT MAP (clk, rst, Multiplier1286Weight, mbRightSHR1286_Input1_1651Output);

    MB_D_FF_Float_1286_1651_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR1286_Input1_1651Output, Multiplier1286WeightOutput);

    InputIEEE_Float_1286_1651: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier1286WeightOutput, flopocoMultiplier1286WeightOutput);

    MB_D_FF_Float_1286_1651_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier1286WeightOutput, flopocoMultiplier1286WeightInput);

    Multiplier_Float_1286: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier1286WeightInput, mb_D_FF1286_1651MultiplierStage2Output, Multiplier1286_Output_1651);

    MBRightSHR_Float_1286_Input2_1651: entity work.MBRightSHR(rtl)
    GENERIC MAP (50, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR1286_Input2_1651Input, mbRightSHR1286_Input2_1651Output);

    MB_D_FF_Float_1286_1651_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR1286_Input2_1651Output, mb_D_FF1286_1651MultiplierStage1Output);

    MB_D_FF_Float_1286_1651_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1286_1651MultiplierStage1Output, mb_D_FF1286_1651MultiplierStage2Output);

    MB_D_FF_Float_Adder16_Input1_365_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier1286_Output_1651, mb_D_FFAdder16_Input1_365_0Output);

    MB_D_FF_Float_365_1652_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder16_Input1_365_0Output, mb_D_FF365_1652AugendStage1Output);

    MB_D_FF_Float_365_1652_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF365_1652AugendStage1Output, mb_D_FF365_1652AugendStage2Output);

    Adder_Float_365: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF365_1652AugendStage2Output, mb_D_FF365_1652AddendStage2Output, Adder365_Output_1652);

    MB_D_FF_Float_Adder16_Input2_365_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier1285_Output_1650, mb_D_FFAdder16_Input2_365_0Output);

    MB_D_FF_Float_365_1652_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder16_Input2_365_0Output, mb_D_FF365_1652AddendStage1Output);

    MB_D_FF_Float_365_1652_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF365_1652AddendStage1Output, mb_D_FF365_1652AddendStage2Output);

    MB_D_FF_Float_Multiplier15_1287_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder365_Output_1652, mb_D_FFMultiplier15_1287_0Output);

    MB_D_FF_Float_1287_1653_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier15_1287_0Output, mb_D_FF1287_1653MultiplierStage1Output);

    MB_D_FF_Float_1287_1653_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1287_1653MultiplierStage1Output, mb_D_FF1287_1653MultiplierStage2Output);

    Multiplier_Float_1287: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF1287_1653MultiplierStage2Output, mb_D_FF1287_1653MultiplicandStage2Output, Multiplier1287_Output_1653);

    MBRightSHR_Float_1287_1653: entity work.MBRightSHR(rtl)
    GENERIC MAP (82, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR1287_1653Input, mbRightSHR1287_1653Output);

    MB_D_FF_Float_1287_1653_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR1287_1653Output, mb_D_FF1287_1653MultiplicandStage1Output);

    MB_D_FF_Float_1287_1653_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1287_1653MultiplicandStage1Output, mb_D_FF1287_1653MultiplicandStage2Output);

    MB_D_FF_Float_Multiplier14_1288_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier1287_Output_1653, mb_D_FFMultiplier14_1288_0Output);

    MB_D_FF_Float_1288_1654_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier14_1288_0Output, mb_D_FF1288_1654MultiplierStage1Output);

    MB_D_FF_Float_1288_1654_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1288_1654MultiplierStage1Output, mb_D_FF1288_1654MultiplierStage2Output);

    Multiplier_Float_1288: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF1288_1654MultiplierStage2Output, flopocoMultiplier1288WeightInput, Multiplier1288_Output_1654);

    MBRightSHR_Float_1288_1654: entity work.MBRightSHR(rtl)
    GENERIC MAP (89, NumberOfBits)
    PORT MAP (clk, rst, Multiplier1288Weight, mbRightSHR1288_1654Output);

    MB_D_FF_Float_1288_1654_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR1288_1654Output, Multiplier1288WeightOutput);

    InputIEEE_Float_1288_1654: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier1288WeightOutput, flopocoMultiplier1288WeightOutput);

    MB_D_FF_Float_1288_1654_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier1288WeightOutput, flopocoMultiplier1288WeightInput);

    MB_D_FF_Float_Multiplier13_1289_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier1288_Output_1654, mb_D_FFMultiplier13_1289_0Output);

    MB_D_FF_Float_1289_1655_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier13_1289_0Output, mb_D_FF1289_1655MultiplierStage1Output);

    MB_D_FF_Float_1289_1655_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1289_1655MultiplierStage1Output, mb_D_FF1289_1655MultiplierStage2Output);

    Multiplier_Float_1289: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF1289_1655MultiplierStage2Output, flopocoMultiplier1289WeightInput, Multiplier1289_Output_1655);

    MBRightSHR_Float_1289_1655: entity work.MBRightSHR(rtl)
    GENERIC MAP (96, NumberOfBits)
    PORT MAP (clk, rst, Multiplier1289Weight, mbRightSHR1289_1655Output);

    MB_D_FF_Float_1289_1655_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR1289_1655Output, Multiplier1289WeightOutput);

    InputIEEE_Float_1289_1655: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier1289WeightOutput, flopocoMultiplier1289WeightOutput);

    MB_D_FF_Float_1289_1655_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier1289WeightOutput, flopocoMultiplier1289WeightInput);

    MBRightSHR_Float_1290_Input11656: entity work.MBRightSHR(rtl)
    GENERIC MAP (50, NumberOfBits)
    PORT MAP (clk, rst, Multiplier1290Weight, mbRightSHR1290_Input1_1656Output);

    MB_D_FF_Float_1290_1656_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR1290_Input1_1656Output, Multiplier1290WeightOutput);

    InputIEEE_Float_1290_1656: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier1290WeightOutput, flopocoMultiplier1290WeightOutput);

    MB_D_FF_Float_1290_1656_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier1290WeightOutput, flopocoMultiplier1290WeightInput);

    Multiplier_Float_1290: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier1290WeightInput, mb_D_FF1290_1656MultiplierStage2Output, Multiplier1290_Output_1656);

    MBRightSHR_Float_1290_Input2_1656: entity work.MBRightSHR(rtl)
    GENERIC MAP (50, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR1290_Input2_1656Input, mbRightSHR1290_Input2_1656Output);

    MB_D_FF_Float_1290_1656_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR1290_Input2_1656Output, mb_D_FF1290_1656MultiplierStage1Output);

    MB_D_FF_Float_1290_1656_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1290_1656MultiplierStage1Output, mb_D_FF1290_1656MultiplierStage2Output);

    MBRightSHR_Float_1291_Input11657: entity work.MBRightSHR(rtl)
    GENERIC MAP (50, NumberOfBits)
    PORT MAP (clk, rst, Multiplier1291Weight, mbRightSHR1291_Input1_1657Output);

    MB_D_FF_Float_1291_1657_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR1291_Input1_1657Output, Multiplier1291WeightOutput);

    InputIEEE_Float_1291_1657: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier1291WeightOutput, flopocoMultiplier1291WeightOutput);

    MB_D_FF_Float_1291_1657_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier1291WeightOutput, flopocoMultiplier1291WeightInput);

    Multiplier_Float_1291: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier1291WeightInput, mb_D_FF1291_1657MultiplierStage2Output, Multiplier1291_Output_1657);

    MBRightSHR_Float_1291_Input2_1657: entity work.MBRightSHR(rtl)
    GENERIC MAP (50, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR1291_Input2_1657Input, mbRightSHR1291_Input2_1657Output);

    MB_D_FF_Float_1291_1657_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR1291_Input2_1657Output, mb_D_FF1291_1657MultiplierStage1Output);

    MB_D_FF_Float_1291_1657_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1291_1657MultiplierStage1Output, mb_D_FF1291_1657MultiplierStage2Output);

    MB_D_FF_Float_Adder16_Input1_366_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier1291_Output_1657, mb_D_FFAdder16_Input1_366_0Output);

    MB_D_FF_Float_366_1658_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder16_Input1_366_0Output, mb_D_FF366_1658AugendStage1Output);

    MB_D_FF_Float_366_1658_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF366_1658AugendStage1Output, mb_D_FF366_1658AugendStage2Output);

    Adder_Float_366: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF366_1658AugendStage2Output, mb_D_FF366_1658AddendStage2Output, Adder366_Output_1658);

    MB_D_FF_Float_Adder16_Input2_366_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier1290_Output_1656, mb_D_FFAdder16_Input2_366_0Output);

    MB_D_FF_Float_366_1658_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder16_Input2_366_0Output, mb_D_FF366_1658AddendStage1Output);

    MB_D_FF_Float_366_1658_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF366_1658AddendStage1Output, mb_D_FF366_1658AddendStage2Output);

    MB_D_FF_Float_Multiplier15_1292_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder366_Output_1658, mb_D_FFMultiplier15_1292_0Output);

    MB_D_FF_Float_1292_1659_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier15_1292_0Output, mb_D_FF1292_1659MultiplierStage1Output);

    MB_D_FF_Float_1292_1659_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1292_1659MultiplierStage1Output, mb_D_FF1292_1659MultiplierStage2Output);

    Multiplier_Float_1292: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF1292_1659MultiplierStage2Output, mb_D_FF1292_1659MultiplicandStage2Output, Multiplier1292_Output_1659);

    MBRightSHR_Float_1292_1659: entity work.MBRightSHR(rtl)
    GENERIC MAP (82, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR1292_1659Input, mbRightSHR1292_1659Output);

    MB_D_FF_Float_1292_1659_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR1292_1659Output, mb_D_FF1292_1659MultiplicandStage1Output);

    MB_D_FF_Float_1292_1659_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1292_1659MultiplicandStage1Output, mb_D_FF1292_1659MultiplicandStage2Output);

    MB_D_FF_Float_Multiplier14_1293_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier1292_Output_1659, mb_D_FFMultiplier14_1293_0Output);

    MB_D_FF_Float_1293_1660_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier14_1293_0Output, mb_D_FF1293_1660MultiplierStage1Output);

    MB_D_FF_Float_1293_1660_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1293_1660MultiplierStage1Output, mb_D_FF1293_1660MultiplierStage2Output);

    Multiplier_Float_1293: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF1293_1660MultiplierStage2Output, flopocoMultiplier1293WeightInput, Multiplier1293_Output_1660);

    MBRightSHR_Float_1293_1660: entity work.MBRightSHR(rtl)
    GENERIC MAP (89, NumberOfBits)
    PORT MAP (clk, rst, Multiplier1293Weight, mbRightSHR1293_1660Output);

    MB_D_FF_Float_1293_1660_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR1293_1660Output, Multiplier1293WeightOutput);

    InputIEEE_Float_1293_1660: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier1293WeightOutput, flopocoMultiplier1293WeightOutput);

    MB_D_FF_Float_1293_1660_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier1293WeightOutput, flopocoMultiplier1293WeightInput);

    MB_D_FF_Float_Multiplier13_1294_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier1293_Output_1660, mb_D_FFMultiplier13_1294_0Output);

    MB_D_FF_Float_1294_1661_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier13_1294_0Output, mb_D_FF1294_1661MultiplierStage1Output);

    MB_D_FF_Float_1294_1661_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1294_1661MultiplierStage1Output, mb_D_FF1294_1661MultiplierStage2Output);

    Multiplier_Float_1294: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF1294_1661MultiplierStage2Output, flopocoMultiplier1294WeightInput, Multiplier1294_Output_1661);

    MBRightSHR_Float_1294_1661: entity work.MBRightSHR(rtl)
    GENERIC MAP (96, NumberOfBits)
    PORT MAP (clk, rst, Multiplier1294Weight, mbRightSHR1294_1661Output);

    MB_D_FF_Float_1294_1661_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR1294_1661Output, Multiplier1294WeightOutput);

    InputIEEE_Float_1294_1661: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier1294WeightOutput, flopocoMultiplier1294WeightOutput);

    MB_D_FF_Float_1294_1661_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier1294WeightOutput, flopocoMultiplier1294WeightInput);

    MB_D_FF_Float_Adder12_Input1_367_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier1294_Output_1661, mb_D_FFAdder12_Input1_367_0Output);

    MB_D_FF_Float_367_1662_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder12_Input1_367_0Output, mb_D_FF367_1662AugendStage1Output);

    MB_D_FF_Float_367_1662_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF367_1662AugendStage1Output, mb_D_FF367_1662AugendStage2Output);

    Adder_Float_367: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF367_1662AugendStage2Output, mb_D_FF367_1662AddendStage2Output, Adder367_Output_1662);

    MB_D_FF_Float_Adder12_Input2_367_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier1289_Output_1655, mb_D_FFAdder12_Input2_367_0Output);

    MB_D_FF_Float_367_1662_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder12_Input2_367_0Output, mb_D_FF367_1662AddendStage1Output);

    MB_D_FF_Float_367_1662_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF367_1662AddendStage1Output, mb_D_FF367_1662AddendStage2Output);

    MB_D_FF_Float_Multiplier11_Input1_1295_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder367_Output_1662, mb_D_FFMultiplier11_Input1_1295_0Output);

    MB_D_FF_Float_1295_1663_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier11_Input1_1295_0Output, mb_D_FF1295_1663MultiplicandStage1Output);

    MB_D_FF_Float_1295_1663_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1295_1663MultiplicandStage1Output, mb_D_FF1295_1663MultiplicandStage2Output);

    Multiplier_Float_1295: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF1295_1663MultiplicandStage2Output, mb_D_FF1295_1663MultiplierStage2Output, Multiplier1295_Output_1663);

    MB_D_FF_Float_Multiplier11_Input2_1295_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier137_Output_171, mb_D_FFMultiplier11_Input2_1295_0Output);

    MB_D_FF_Float_1295_1663_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier11_Input2_1295_0Output, mb_D_FF1295_1663MultiplierStage1Output);

    MB_D_FF_Float_1295_1663_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1295_1663MultiplierStage1Output, mb_D_FF1295_1663MultiplierStage2Output);

    MBRightSHR_Float_1329_Input11708: entity work.MBRightSHR(rtl)
    GENERIC MAP (50, NumberOfBits)
    PORT MAP (clk, rst, Multiplier1329Weight, mbRightSHR1329_Input1_1708Output);

    MB_D_FF_Float_1329_1708_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR1329_Input1_1708Output, Multiplier1329WeightOutput);

    InputIEEE_Float_1329_1708: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier1329WeightOutput, flopocoMultiplier1329WeightOutput);

    MB_D_FF_Float_1329_1708_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier1329WeightOutput, flopocoMultiplier1329WeightInput);

    Multiplier_Float_1329: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier1329WeightInput, mb_D_FF1329_1708MultiplierStage2Output, Multiplier1329_Output_1708);

    MBRightSHR_Float_1329_Input2_1708: entity work.MBRightSHR(rtl)
    GENERIC MAP (50, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR1329_Input2_1708Input, mbRightSHR1329_Input2_1708Output);

    MB_D_FF_Float_1329_1708_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR1329_Input2_1708Output, mb_D_FF1329_1708MultiplierStage1Output);

    MB_D_FF_Float_1329_1708_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1329_1708MultiplierStage1Output, mb_D_FF1329_1708MultiplierStage2Output);

    MBRightSHR_Float_1330_Input11709: entity work.MBRightSHR(rtl)
    GENERIC MAP (50, NumberOfBits)
    PORT MAP (clk, rst, Multiplier1330Weight, mbRightSHR1330_Input1_1709Output);

    MB_D_FF_Float_1330_1709_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR1330_Input1_1709Output, Multiplier1330WeightOutput);

    InputIEEE_Float_1330_1709: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier1330WeightOutput, flopocoMultiplier1330WeightOutput);

    MB_D_FF_Float_1330_1709_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier1330WeightOutput, flopocoMultiplier1330WeightInput);

    Multiplier_Float_1330: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier1330WeightInput, mb_D_FF1330_1709MultiplierStage2Output, Multiplier1330_Output_1709);

    MBRightSHR_Float_1330_Input2_1709: entity work.MBRightSHR(rtl)
    GENERIC MAP (50, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR1330_Input2_1709Input, mbRightSHR1330_Input2_1709Output);

    MB_D_FF_Float_1330_1709_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR1330_Input2_1709Output, mb_D_FF1330_1709MultiplierStage1Output);

    MB_D_FF_Float_1330_1709_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1330_1709MultiplierStage1Output, mb_D_FF1330_1709MultiplierStage2Output);

    MB_D_FF_Float_Adder16_Input1_379_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier1330_Output_1709, mb_D_FFAdder16_Input1_379_0Output);

    MB_D_FF_Float_379_1710_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder16_Input1_379_0Output, mb_D_FF379_1710AugendStage1Output);

    MB_D_FF_Float_379_1710_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF379_1710AugendStage1Output, mb_D_FF379_1710AugendStage2Output);

    Adder_Float_379: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF379_1710AugendStage2Output, mb_D_FF379_1710AddendStage2Output, Adder379_Output_1710);

    MB_D_FF_Float_Adder16_Input2_379_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier1329_Output_1708, mb_D_FFAdder16_Input2_379_0Output);

    MB_D_FF_Float_379_1710_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder16_Input2_379_0Output, mb_D_FF379_1710AddendStage1Output);

    MB_D_FF_Float_379_1710_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF379_1710AddendStage1Output, mb_D_FF379_1710AddendStage2Output);

    MB_D_FF_Float_Multiplier15_1331_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder379_Output_1710, mb_D_FFMultiplier15_1331_0Output);

    MB_D_FF_Float_1331_1711_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier15_1331_0Output, mb_D_FF1331_1711MultiplierStage1Output);

    MB_D_FF_Float_1331_1711_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1331_1711MultiplierStage1Output, mb_D_FF1331_1711MultiplierStage2Output);

    Multiplier_Float_1331: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF1331_1711MultiplierStage2Output, mb_D_FF1331_1711MultiplicandStage2Output, Multiplier1331_Output_1711);

    MBRightSHR_Float_1331_1711: entity work.MBRightSHR(rtl)
    GENERIC MAP (82, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR1331_1711Input, mbRightSHR1331_1711Output);

    MB_D_FF_Float_1331_1711_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR1331_1711Output, mb_D_FF1331_1711MultiplicandStage1Output);

    MB_D_FF_Float_1331_1711_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1331_1711MultiplicandStage1Output, mb_D_FF1331_1711MultiplicandStage2Output);

    MB_D_FF_Float_Multiplier14_1332_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier1331_Output_1711, mb_D_FFMultiplier14_1332_0Output);

    MB_D_FF_Float_1332_1712_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier14_1332_0Output, mb_D_FF1332_1712MultiplierStage1Output);

    MB_D_FF_Float_1332_1712_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1332_1712MultiplierStage1Output, mb_D_FF1332_1712MultiplierStage2Output);

    Multiplier_Float_1332: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF1332_1712MultiplierStage2Output, flopocoMultiplier1332WeightInput, Multiplier1332_Output_1712);

    MBRightSHR_Float_1332_1712: entity work.MBRightSHR(rtl)
    GENERIC MAP (89, NumberOfBits)
    PORT MAP (clk, rst, Multiplier1332Weight, mbRightSHR1332_1712Output);

    MB_D_FF_Float_1332_1712_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR1332_1712Output, Multiplier1332WeightOutput);

    InputIEEE_Float_1332_1712: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier1332WeightOutput, flopocoMultiplier1332WeightOutput);

    MB_D_FF_Float_1332_1712_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier1332WeightOutput, flopocoMultiplier1332WeightInput);

    MB_D_FF_Float_Multiplier13_1333_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier1332_Output_1712, mb_D_FFMultiplier13_1333_0Output);

    MB_D_FF_Float_1333_1713_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier13_1333_0Output, mb_D_FF1333_1713MultiplierStage1Output);

    MB_D_FF_Float_1333_1713_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1333_1713MultiplierStage1Output, mb_D_FF1333_1713MultiplierStage2Output);

    Multiplier_Float_1333: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF1333_1713MultiplierStage2Output, flopocoMultiplier1333WeightInput, Multiplier1333_Output_1713);

    MBRightSHR_Float_1333_1713: entity work.MBRightSHR(rtl)
    GENERIC MAP (96, NumberOfBits)
    PORT MAP (clk, rst, Multiplier1333Weight, mbRightSHR1333_1713Output);

    MB_D_FF_Float_1333_1713_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR1333_1713Output, Multiplier1333WeightOutput);

    InputIEEE_Float_1333_1713: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier1333WeightOutput, flopocoMultiplier1333WeightOutput);

    MB_D_FF_Float_1333_1713_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier1333WeightOutput, flopocoMultiplier1333WeightInput);

    MBRightSHR_Float_1334_Input11714: entity work.MBRightSHR(rtl)
    GENERIC MAP (50, NumberOfBits)
    PORT MAP (clk, rst, Multiplier1334Weight, mbRightSHR1334_Input1_1714Output);

    MB_D_FF_Float_1334_1714_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR1334_Input1_1714Output, Multiplier1334WeightOutput);

    InputIEEE_Float_1334_1714: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier1334WeightOutput, flopocoMultiplier1334WeightOutput);

    MB_D_FF_Float_1334_1714_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier1334WeightOutput, flopocoMultiplier1334WeightInput);

    Multiplier_Float_1334: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier1334WeightInput, mb_D_FF1334_1714MultiplierStage2Output, Multiplier1334_Output_1714);

    MBRightSHR_Float_1334_Input2_1714: entity work.MBRightSHR(rtl)
    GENERIC MAP (50, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR1334_Input2_1714Input, mbRightSHR1334_Input2_1714Output);

    MB_D_FF_Float_1334_1714_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR1334_Input2_1714Output, mb_D_FF1334_1714MultiplierStage1Output);

    MB_D_FF_Float_1334_1714_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1334_1714MultiplierStage1Output, mb_D_FF1334_1714MultiplierStage2Output);

    MBRightSHR_Float_1335_Input11715: entity work.MBRightSHR(rtl)
    GENERIC MAP (50, NumberOfBits)
    PORT MAP (clk, rst, Multiplier1335Weight, mbRightSHR1335_Input1_1715Output);

    MB_D_FF_Float_1335_1715_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR1335_Input1_1715Output, Multiplier1335WeightOutput);

    InputIEEE_Float_1335_1715: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier1335WeightOutput, flopocoMultiplier1335WeightOutput);

    MB_D_FF_Float_1335_1715_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier1335WeightOutput, flopocoMultiplier1335WeightInput);

    Multiplier_Float_1335: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier1335WeightInput, mb_D_FF1335_1715MultiplierStage2Output, Multiplier1335_Output_1715);

    MBRightSHR_Float_1335_Input2_1715: entity work.MBRightSHR(rtl)
    GENERIC MAP (50, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR1335_Input2_1715Input, mbRightSHR1335_Input2_1715Output);

    MB_D_FF_Float_1335_1715_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR1335_Input2_1715Output, mb_D_FF1335_1715MultiplierStage1Output);

    MB_D_FF_Float_1335_1715_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1335_1715MultiplierStage1Output, mb_D_FF1335_1715MultiplierStage2Output);

    MB_D_FF_Float_Adder16_Input1_380_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier1335_Output_1715, mb_D_FFAdder16_Input1_380_0Output);

    MB_D_FF_Float_380_1716_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder16_Input1_380_0Output, mb_D_FF380_1716AugendStage1Output);

    MB_D_FF_Float_380_1716_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF380_1716AugendStage1Output, mb_D_FF380_1716AugendStage2Output);

    Adder_Float_380: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF380_1716AugendStage2Output, mb_D_FF380_1716AddendStage2Output, Adder380_Output_1716);

    MB_D_FF_Float_Adder16_Input2_380_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier1334_Output_1714, mb_D_FFAdder16_Input2_380_0Output);

    MB_D_FF_Float_380_1716_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder16_Input2_380_0Output, mb_D_FF380_1716AddendStage1Output);

    MB_D_FF_Float_380_1716_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF380_1716AddendStage1Output, mb_D_FF380_1716AddendStage2Output);

    MB_D_FF_Float_Multiplier15_1336_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder380_Output_1716, mb_D_FFMultiplier15_1336_0Output);

    MB_D_FF_Float_1336_1717_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier15_1336_0Output, mb_D_FF1336_1717MultiplierStage1Output);

    MB_D_FF_Float_1336_1717_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1336_1717MultiplierStage1Output, mb_D_FF1336_1717MultiplierStage2Output);

    Multiplier_Float_1336: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF1336_1717MultiplierStage2Output, mb_D_FF1336_1717MultiplicandStage2Output, Multiplier1336_Output_1717);

    MBRightSHR_Float_1336_1717: entity work.MBRightSHR(rtl)
    GENERIC MAP (82, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR1336_1717Input, mbRightSHR1336_1717Output);

    MB_D_FF_Float_1336_1717_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR1336_1717Output, mb_D_FF1336_1717MultiplicandStage1Output);

    MB_D_FF_Float_1336_1717_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1336_1717MultiplicandStage1Output, mb_D_FF1336_1717MultiplicandStage2Output);

    MB_D_FF_Float_Multiplier14_1337_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier1336_Output_1717, mb_D_FFMultiplier14_1337_0Output);

    MB_D_FF_Float_1337_1718_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier14_1337_0Output, mb_D_FF1337_1718MultiplierStage1Output);

    MB_D_FF_Float_1337_1718_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1337_1718MultiplierStage1Output, mb_D_FF1337_1718MultiplierStage2Output);

    Multiplier_Float_1337: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF1337_1718MultiplierStage2Output, flopocoMultiplier1337WeightInput, Multiplier1337_Output_1718);

    MBRightSHR_Float_1337_1718: entity work.MBRightSHR(rtl)
    GENERIC MAP (89, NumberOfBits)
    PORT MAP (clk, rst, Multiplier1337Weight, mbRightSHR1337_1718Output);

    MB_D_FF_Float_1337_1718_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR1337_1718Output, Multiplier1337WeightOutput);

    InputIEEE_Float_1337_1718: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier1337WeightOutput, flopocoMultiplier1337WeightOutput);

    MB_D_FF_Float_1337_1718_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier1337WeightOutput, flopocoMultiplier1337WeightInput);

    MB_D_FF_Float_Multiplier13_1338_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier1337_Output_1718, mb_D_FFMultiplier13_1338_0Output);

    MB_D_FF_Float_1338_1719_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier13_1338_0Output, mb_D_FF1338_1719MultiplierStage1Output);

    MB_D_FF_Float_1338_1719_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1338_1719MultiplierStage1Output, mb_D_FF1338_1719MultiplierStage2Output);

    Multiplier_Float_1338: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF1338_1719MultiplierStage2Output, flopocoMultiplier1338WeightInput, Multiplier1338_Output_1719);

    MBRightSHR_Float_1338_1719: entity work.MBRightSHR(rtl)
    GENERIC MAP (96, NumberOfBits)
    PORT MAP (clk, rst, Multiplier1338Weight, mbRightSHR1338_1719Output);

    MB_D_FF_Float_1338_1719_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR1338_1719Output, Multiplier1338WeightOutput);

    InputIEEE_Float_1338_1719: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier1338WeightOutput, flopocoMultiplier1338WeightOutput);

    MB_D_FF_Float_1338_1719_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier1338WeightOutput, flopocoMultiplier1338WeightInput);

    MB_D_FF_Float_Adder12_Input1_381_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier1338_Output_1719, mb_D_FFAdder12_Input1_381_0Output);

    MB_D_FF_Float_381_1720_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder12_Input1_381_0Output, mb_D_FF381_1720AugendStage1Output);

    MB_D_FF_Float_381_1720_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF381_1720AugendStage1Output, mb_D_FF381_1720AugendStage2Output);

    Adder_Float_381: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF381_1720AugendStage2Output, mb_D_FF381_1720AddendStage2Output, Adder381_Output_1720);

    MB_D_FF_Float_Adder12_Input2_381_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier1333_Output_1713, mb_D_FFAdder12_Input2_381_0Output);

    MB_D_FF_Float_381_1720_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder12_Input2_381_0Output, mb_D_FF381_1720AddendStage1Output);

    MB_D_FF_Float_381_1720_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF381_1720AddendStage1Output, mb_D_FF381_1720AddendStage2Output);

    MB_D_FF_Float_Multiplier11_Input1_1339_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder381_Output_1720, mb_D_FFMultiplier11_Input1_1339_0Output);

    MB_D_FF_Float_1339_1721_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier11_Input1_1339_0Output, mb_D_FF1339_1721MultiplicandStage1Output);

    MB_D_FF_Float_1339_1721_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1339_1721MultiplicandStage1Output, mb_D_FF1339_1721MultiplicandStage2Output);

    Multiplier_Float_1339: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF1339_1721MultiplicandStage2Output, mb_D_FF1339_1721MultiplierStage2Output, Multiplier1339_Output_1721);

    MB_D_FF_Float_Multiplier11_Input2_1339_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier181_Output_229, mb_D_FFMultiplier11_Input2_1339_0Output);

    MB_D_FF_Float_1339_1721_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier11_Input2_1339_0Output, mb_D_FF1339_1721MultiplierStage1Output);

    MB_D_FF_Float_1339_1721_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1339_1721MultiplierStage1Output, mb_D_FF1339_1721MultiplierStage2Output);

    MB_D_FF_Float_Adder10_Input1_382_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier1339_Output_1721, mb_D_FFAdder10_Input1_382_0Output);

    MB_D_FF_Float_382_1722_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder10_Input1_382_0Output, mb_D_FF382_1722AugendStage1Output);

    MB_D_FF_Float_382_1722_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF382_1722AugendStage1Output, mb_D_FF382_1722AugendStage2Output);

    Adder_Float_382: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF382_1722AugendStage2Output, mb_D_FF382_1722AddendStage2Output, Adder382_Output_1722);

    MB_D_FF_Float_Adder10_Input2_382_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier1295_Output_1663, mb_D_FFAdder10_Input2_382_0Output);

    MB_D_FF_Float_382_1722_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder10_Input2_382_0Output, mb_D_FF382_1722AddendStage1Output);

    MB_D_FF_Float_382_1722_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF382_1722AddendStage1Output, mb_D_FF382_1722AddendStage2Output);

    MB_D_FF_Float_Multiplier9_1340_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder382_Output_1722, mb_D_FFMultiplier9_1340_0Output);

    MB_D_FF_Float_1340_1723_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier9_1340_0Output, mb_D_FF1340_1723MultiplierStage1Output);

    MB_D_FF_Float_1340_1723_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1340_1723MultiplierStage1Output, mb_D_FF1340_1723MultiplierStage2Output);

    Multiplier_Float_1340: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF1340_1723MultiplierStage2Output, mb_D_FF1340_1723MultiplicandStage2Output, Multiplier1340_Output_1723);

    MBRightSHR_Float_1340_1723: entity work.MBRightSHR(rtl)
    GENERIC MAP (160, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR1340_1723Input, mbRightSHR1340_1723Output);

    MB_D_FF_Float_1340_1723_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR1340_1723Output, mb_D_FF1340_1723MultiplicandStage1Output);

    MB_D_FF_Float_1340_1723_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1340_1723MultiplicandStage1Output, mb_D_FF1340_1723MultiplicandStage2Output);

    MB_D_FF_Float_Multiplier8_1341_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier1340_Output_1723, mb_D_FFMultiplier8_1341_0Output);

    MB_D_FF_Float_1341_1724_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier8_1341_0Output, mb_D_FF1341_1724MultiplierStage1Output);

    MB_D_FF_Float_1341_1724_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1341_1724MultiplierStage1Output, mb_D_FF1341_1724MultiplierStage2Output);

    Multiplier_Float_1341: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF1341_1724MultiplierStage2Output, flopocoMultiplier1341WeightInput, Multiplier1341_Output_1724);

    MBRightSHR_Float_1341_1724: entity work.MBRightSHR(rtl)
    GENERIC MAP (167, NumberOfBits)
    PORT MAP (clk, rst, Multiplier1341Weight, mbRightSHR1341_1724Output);

    MB_D_FF_Float_1341_1724_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR1341_1724Output, Multiplier1341WeightOutput);

    InputIEEE_Float_1341_1724: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier1341WeightOutput, flopocoMultiplier1341WeightOutput);

    MB_D_FF_Float_1341_1724_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier1341WeightOutput, flopocoMultiplier1341WeightInput);

    MB_D_FF_Float_Multiplier14_1378_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier1287_Output_1653, mb_D_FFMultiplier14_1378_0Output);

    MB_D_FF_Float_1378_1773_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier14_1378_0Output, mb_D_FF1378_1773MultiplierStage1Output);

    MB_D_FF_Float_1378_1773_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1378_1773MultiplierStage1Output, mb_D_FF1378_1773MultiplierStage2Output);

    Multiplier_Float_1378: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF1378_1773MultiplierStage2Output, flopocoMultiplier1378WeightInput, Multiplier1378_Output_1773);

    MBRightSHR_Float_1378_1773: entity work.MBRightSHR(rtl)
    GENERIC MAP (89, NumberOfBits)
    PORT MAP (clk, rst, Multiplier1378Weight, mbRightSHR1378_1773Output);

    MB_D_FF_Float_1378_1773_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR1378_1773Output, Multiplier1378WeightOutput);

    InputIEEE_Float_1378_1773: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier1378WeightOutput, flopocoMultiplier1378WeightOutput);

    MB_D_FF_Float_1378_1773_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier1378WeightOutput, flopocoMultiplier1378WeightInput);

    MB_D_FF_Float_Multiplier13_1379_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier1378_Output_1773, mb_D_FFMultiplier13_1379_0Output);

    MB_D_FF_Float_1379_1774_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier13_1379_0Output, mb_D_FF1379_1774MultiplierStage1Output);

    MB_D_FF_Float_1379_1774_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1379_1774MultiplierStage1Output, mb_D_FF1379_1774MultiplierStage2Output);

    Multiplier_Float_1379: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF1379_1774MultiplierStage2Output, flopocoMultiplier1379WeightInput, Multiplier1379_Output_1774);

    MBRightSHR_Float_1379_1774: entity work.MBRightSHR(rtl)
    GENERIC MAP (96, NumberOfBits)
    PORT MAP (clk, rst, Multiplier1379Weight, mbRightSHR1379_1774Output);

    MB_D_FF_Float_1379_1774_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR1379_1774Output, Multiplier1379WeightOutput);

    InputIEEE_Float_1379_1774: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier1379WeightOutput, flopocoMultiplier1379WeightOutput);

    MB_D_FF_Float_1379_1774_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier1379WeightOutput, flopocoMultiplier1379WeightInput);

    MB_D_FF_Float_Multiplier14_1383_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier1292_Output_1659, mb_D_FFMultiplier14_1383_0Output);

    MB_D_FF_Float_1383_1779_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier14_1383_0Output, mb_D_FF1383_1779MultiplierStage1Output);

    MB_D_FF_Float_1383_1779_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1383_1779MultiplierStage1Output, mb_D_FF1383_1779MultiplierStage2Output);

    Multiplier_Float_1383: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF1383_1779MultiplierStage2Output, flopocoMultiplier1383WeightInput, Multiplier1383_Output_1779);

    MBRightSHR_Float_1383_1779: entity work.MBRightSHR(rtl)
    GENERIC MAP (89, NumberOfBits)
    PORT MAP (clk, rst, Multiplier1383Weight, mbRightSHR1383_1779Output);

    MB_D_FF_Float_1383_1779_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR1383_1779Output, Multiplier1383WeightOutput);

    InputIEEE_Float_1383_1779: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier1383WeightOutput, flopocoMultiplier1383WeightOutput);

    MB_D_FF_Float_1383_1779_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier1383WeightOutput, flopocoMultiplier1383WeightInput);

    MB_D_FF_Float_Multiplier13_1384_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier1383_Output_1779, mb_D_FFMultiplier13_1384_0Output);

    MB_D_FF_Float_1384_1780_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier13_1384_0Output, mb_D_FF1384_1780MultiplierStage1Output);

    MB_D_FF_Float_1384_1780_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1384_1780MultiplierStage1Output, mb_D_FF1384_1780MultiplierStage2Output);

    Multiplier_Float_1384: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF1384_1780MultiplierStage2Output, flopocoMultiplier1384WeightInput, Multiplier1384_Output_1780);

    MBRightSHR_Float_1384_1780: entity work.MBRightSHR(rtl)
    GENERIC MAP (96, NumberOfBits)
    PORT MAP (clk, rst, Multiplier1384Weight, mbRightSHR1384_1780Output);

    MB_D_FF_Float_1384_1780_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR1384_1780Output, Multiplier1384WeightOutput);

    InputIEEE_Float_1384_1780: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier1384WeightOutput, flopocoMultiplier1384WeightOutput);

    MB_D_FF_Float_1384_1780_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier1384WeightOutput, flopocoMultiplier1384WeightInput);

    MB_D_FF_Float_Adder12_Input1_396_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier1384_Output_1780, mb_D_FFAdder12_Input1_396_0Output);

    MB_D_FF_Float_396_1781_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder12_Input1_396_0Output, mb_D_FF396_1781AugendStage1Output);

    MB_D_FF_Float_396_1781_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF396_1781AugendStage1Output, mb_D_FF396_1781AugendStage2Output);

    Adder_Float_396: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF396_1781AugendStage2Output, mb_D_FF396_1781AddendStage2Output, Adder396_Output_1781);

    MB_D_FF_Float_Adder12_Input2_396_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier1379_Output_1774, mb_D_FFAdder12_Input2_396_0Output);

    MB_D_FF_Float_396_1781_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder12_Input2_396_0Output, mb_D_FF396_1781AddendStage1Output);

    MB_D_FF_Float_396_1781_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF396_1781AddendStage1Output, mb_D_FF396_1781AddendStage2Output);

    MB_D_FF_Float_Multiplier11_Input1_1385_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder396_Output_1781, mb_D_FFMultiplier11_Input1_1385_0Output);

    MB_D_FF_Float_1385_1782_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier11_Input1_1385_0Output, mb_D_FF1385_1782MultiplicandStage1Output);

    MB_D_FF_Float_1385_1782_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1385_1782MultiplicandStage1Output, mb_D_FF1385_1782MultiplicandStage2Output);

    Multiplier_Float_1385: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF1385_1782MultiplicandStage2Output, mb_D_FF1385_1782MultiplierStage2Output, Multiplier1385_Output_1782);

    MB_D_FF_Float_Multiplier11_Input2_1385_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier227_Output_290, mb_D_FFMultiplier11_Input2_1385_0Output);

    MB_D_FF_Float_1385_1782_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier11_Input2_1385_0Output, mb_D_FF1385_1782MultiplierStage1Output);

    MB_D_FF_Float_1385_1782_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1385_1782MultiplierStage1Output, mb_D_FF1385_1782MultiplierStage2Output);

    MB_D_FF_Float_Multiplier14_1422_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier1331_Output_1711, mb_D_FFMultiplier14_1422_0Output);

    MB_D_FF_Float_1422_1831_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier14_1422_0Output, mb_D_FF1422_1831MultiplierStage1Output);

    MB_D_FF_Float_1422_1831_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1422_1831MultiplierStage1Output, mb_D_FF1422_1831MultiplierStage2Output);

    Multiplier_Float_1422: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF1422_1831MultiplierStage2Output, flopocoMultiplier1422WeightInput, Multiplier1422_Output_1831);

    MBRightSHR_Float_1422_1831: entity work.MBRightSHR(rtl)
    GENERIC MAP (89, NumberOfBits)
    PORT MAP (clk, rst, Multiplier1422Weight, mbRightSHR1422_1831Output);

    MB_D_FF_Float_1422_1831_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR1422_1831Output, Multiplier1422WeightOutput);

    InputIEEE_Float_1422_1831: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier1422WeightOutput, flopocoMultiplier1422WeightOutput);

    MB_D_FF_Float_1422_1831_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier1422WeightOutput, flopocoMultiplier1422WeightInput);

    MB_D_FF_Float_Multiplier13_1423_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier1422_Output_1831, mb_D_FFMultiplier13_1423_0Output);

    MB_D_FF_Float_1423_1832_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier13_1423_0Output, mb_D_FF1423_1832MultiplierStage1Output);

    MB_D_FF_Float_1423_1832_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1423_1832MultiplierStage1Output, mb_D_FF1423_1832MultiplierStage2Output);

    Multiplier_Float_1423: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF1423_1832MultiplierStage2Output, flopocoMultiplier1423WeightInput, Multiplier1423_Output_1832);

    MBRightSHR_Float_1423_1832: entity work.MBRightSHR(rtl)
    GENERIC MAP (96, NumberOfBits)
    PORT MAP (clk, rst, Multiplier1423Weight, mbRightSHR1423_1832Output);

    MB_D_FF_Float_1423_1832_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR1423_1832Output, Multiplier1423WeightOutput);

    InputIEEE_Float_1423_1832: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier1423WeightOutput, flopocoMultiplier1423WeightOutput);

    MB_D_FF_Float_1423_1832_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier1423WeightOutput, flopocoMultiplier1423WeightInput);

    MB_D_FF_Float_Multiplier14_1427_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier1336_Output_1717, mb_D_FFMultiplier14_1427_0Output);

    MB_D_FF_Float_1427_1837_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier14_1427_0Output, mb_D_FF1427_1837MultiplierStage1Output);

    MB_D_FF_Float_1427_1837_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1427_1837MultiplierStage1Output, mb_D_FF1427_1837MultiplierStage2Output);

    Multiplier_Float_1427: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF1427_1837MultiplierStage2Output, flopocoMultiplier1427WeightInput, Multiplier1427_Output_1837);

    MBRightSHR_Float_1427_1837: entity work.MBRightSHR(rtl)
    GENERIC MAP (89, NumberOfBits)
    PORT MAP (clk, rst, Multiplier1427Weight, mbRightSHR1427_1837Output);

    MB_D_FF_Float_1427_1837_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR1427_1837Output, Multiplier1427WeightOutput);

    InputIEEE_Float_1427_1837: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier1427WeightOutput, flopocoMultiplier1427WeightOutput);

    MB_D_FF_Float_1427_1837_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier1427WeightOutput, flopocoMultiplier1427WeightInput);

    MB_D_FF_Float_Multiplier13_1428_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier1427_Output_1837, mb_D_FFMultiplier13_1428_0Output);

    MB_D_FF_Float_1428_1838_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier13_1428_0Output, mb_D_FF1428_1838MultiplierStage1Output);

    MB_D_FF_Float_1428_1838_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1428_1838MultiplierStage1Output, mb_D_FF1428_1838MultiplierStage2Output);

    Multiplier_Float_1428: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF1428_1838MultiplierStage2Output, flopocoMultiplier1428WeightInput, Multiplier1428_Output_1838);

    MBRightSHR_Float_1428_1838: entity work.MBRightSHR(rtl)
    GENERIC MAP (96, NumberOfBits)
    PORT MAP (clk, rst, Multiplier1428Weight, mbRightSHR1428_1838Output);

    MB_D_FF_Float_1428_1838_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR1428_1838Output, Multiplier1428WeightOutput);

    InputIEEE_Float_1428_1838: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier1428WeightOutput, flopocoMultiplier1428WeightOutput);

    MB_D_FF_Float_1428_1838_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier1428WeightOutput, flopocoMultiplier1428WeightInput);

    MB_D_FF_Float_Adder12_Input1_410_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier1428_Output_1838, mb_D_FFAdder12_Input1_410_0Output);

    MB_D_FF_Float_410_1839_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder12_Input1_410_0Output, mb_D_FF410_1839AugendStage1Output);

    MB_D_FF_Float_410_1839_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF410_1839AugendStage1Output, mb_D_FF410_1839AugendStage2Output);

    Adder_Float_410: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF410_1839AugendStage2Output, mb_D_FF410_1839AddendStage2Output, Adder410_Output_1839);

    MB_D_FF_Float_Adder12_Input2_410_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier1423_Output_1832, mb_D_FFAdder12_Input2_410_0Output);

    MB_D_FF_Float_410_1839_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder12_Input2_410_0Output, mb_D_FF410_1839AddendStage1Output);

    MB_D_FF_Float_410_1839_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF410_1839AddendStage1Output, mb_D_FF410_1839AddendStage2Output);

    MB_D_FF_Float_Multiplier11_Input1_1429_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder410_Output_1839, mb_D_FFMultiplier11_Input1_1429_0Output);

    MB_D_FF_Float_1429_1840_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier11_Input1_1429_0Output, mb_D_FF1429_1840MultiplicandStage1Output);

    MB_D_FF_Float_1429_1840_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1429_1840MultiplicandStage1Output, mb_D_FF1429_1840MultiplicandStage2Output);

    Multiplier_Float_1429: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF1429_1840MultiplicandStage2Output, mb_D_FF1429_1840MultiplierStage2Output, Multiplier1429_Output_1840);

    MB_D_FF_Float_Multiplier11_Input2_1429_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier271_Output_348, mb_D_FFMultiplier11_Input2_1429_0Output);

    MB_D_FF_Float_1429_1840_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier11_Input2_1429_0Output, mb_D_FF1429_1840MultiplierStage1Output);

    MB_D_FF_Float_1429_1840_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1429_1840MultiplierStage1Output, mb_D_FF1429_1840MultiplierStage2Output);

    MB_D_FF_Float_Adder10_Input1_411_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier1429_Output_1840, mb_D_FFAdder10_Input1_411_0Output);

    MB_D_FF_Float_411_1841_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder10_Input1_411_0Output, mb_D_FF411_1841AugendStage1Output);

    MB_D_FF_Float_411_1841_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF411_1841AugendStage1Output, mb_D_FF411_1841AugendStage2Output);

    Adder_Float_411: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF411_1841AugendStage2Output, mb_D_FF411_1841AddendStage2Output, Adder411_Output_1841);

    MB_D_FF_Float_Adder10_Input2_411_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier1385_Output_1782, mb_D_FFAdder10_Input2_411_0Output);

    MB_D_FF_Float_411_1841_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder10_Input2_411_0Output, mb_D_FF411_1841AddendStage1Output);

    MB_D_FF_Float_411_1841_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF411_1841AddendStage1Output, mb_D_FF411_1841AddendStage2Output);

    MB_D_FF_Float_Multiplier9_1430_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder411_Output_1841, mb_D_FFMultiplier9_1430_0Output);

    MB_D_FF_Float_1430_1842_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier9_1430_0Output, mb_D_FF1430_1842MultiplierStage1Output);

    MB_D_FF_Float_1430_1842_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1430_1842MultiplierStage1Output, mb_D_FF1430_1842MultiplierStage2Output);

    Multiplier_Float_1430: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF1430_1842MultiplierStage2Output, mb_D_FF1430_1842MultiplicandStage2Output, Multiplier1430_Output_1842);

    MBRightSHR_Float_1430_1842: entity work.MBRightSHR(rtl)
    GENERIC MAP (160, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR1430_1842Input, mbRightSHR1430_1842Output);

    MB_D_FF_Float_1430_1842_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR1430_1842Output, mb_D_FF1430_1842MultiplicandStage1Output);

    MB_D_FF_Float_1430_1842_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1430_1842MultiplicandStage1Output, mb_D_FF1430_1842MultiplicandStage2Output);

    MB_D_FF_Float_Multiplier8_1431_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier1430_Output_1842, mb_D_FFMultiplier8_1431_0Output);

    MB_D_FF_Float_1431_1843_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier8_1431_0Output, mb_D_FF1431_1843MultiplierStage1Output);

    MB_D_FF_Float_1431_1843_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1431_1843MultiplierStage1Output, mb_D_FF1431_1843MultiplierStage2Output);

    Multiplier_Float_1431: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF1431_1843MultiplierStage2Output, flopocoMultiplier1431WeightInput, Multiplier1431_Output_1843);

    MBRightSHR_Float_1431_1843: entity work.MBRightSHR(rtl)
    GENERIC MAP (167, NumberOfBits)
    PORT MAP (clk, rst, Multiplier1431Weight, mbRightSHR1431_1843Output);

    MB_D_FF_Float_1431_1843_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR1431_1843Output, Multiplier1431WeightOutput);

    InputIEEE_Float_1431_1843: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier1431WeightOutput, flopocoMultiplier1431WeightOutput);

    MB_D_FF_Float_1431_1843_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier1431WeightOutput, flopocoMultiplier1431WeightInput);

    MB_D_FF_Float_Adder7_Input1_412_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier1431_Output_1843, mb_D_FFAdder7_Input1_412_0Output);

    MB_D_FF_Float_412_1844_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder7_Input1_412_0Output, mb_D_FF412_1844AugendStage1Output);

    MB_D_FF_Float_412_1844_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF412_1844AugendStage1Output, mb_D_FF412_1844AugendStage2Output);

    Adder_Float_412: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF412_1844AugendStage2Output, mb_D_FF412_1844AddendStage2Output, Adder412_Output_1844);

    MB_D_FF_Float_Adder7_Input2_412_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier1341_Output_1724, mb_D_FFAdder7_Input2_412_0Output);

    MB_D_FF_Float_412_1844_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder7_Input2_412_0Output, mb_D_FF412_1844AddendStage1Output);

    MB_D_FF_Float_412_1844_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF412_1844AddendStage1Output, mb_D_FF412_1844AddendStage2Output);

    MB_D_FF_Float_Multiplier6_Input1_1432_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder412_Output_1844, mb_D_FFMultiplier6_Input1_1432_0Output);

    MB_D_FF_Float_1432_1845_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier6_Input1_1432_0Output, mb_D_FF1432_1845MultiplicandStage1Output);

    MB_D_FF_Float_1432_1845_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1432_1845MultiplicandStage1Output, mb_D_FF1432_1845MultiplicandStage2Output);

    Multiplier_Float_1432: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF1432_1845MultiplicandStage2Output, mb_D_FF1432_1845MultiplierStage2Output, Multiplier1432_Output_1845);

    MB_D_FF_Float_Multiplier6_Input2_1432_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier1251_Output_1605, mb_D_FFMultiplier6_Input2_1432_0Output);

    MB_D_FF_Float_1432_1845_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier6_Input2_1432_0Output, mb_D_FF1432_1845MultiplierStage1Output);

    MB_D_FF_Float_1432_1845_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1432_1845MultiplierStage1Output, mb_D_FF1432_1845MultiplierStage2Output);

    MB_D_FF_Float_Multiplier9_1484_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier336_Output_429, mb_D_FFMultiplier9_1484_0Output);

    MB_D_FF_Float_1484_1908_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier9_1484_0Output, mb_D_FF1484_1908MultiplierStage1Output);

    MB_D_FF_Float_1484_1908_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1484_1908MultiplierStage1Output, mb_D_FF1484_1908MultiplierStage2Output);

    Multiplier_Float_1484: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF1484_1908MultiplierStage2Output, flopocoMultiplier1484WeightInput, Multiplier1484_Output_1908);

    MBRightSHR_Float_1484_1908: entity work.MBRightSHR(rtl)
    GENERIC MAP (160, NumberOfBits)
    PORT MAP (clk, rst, Multiplier1484Weight, mbRightSHR1484_1908Output);

    MB_D_FF_Float_1484_1908_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR1484_1908Output, Multiplier1484WeightOutput);

    InputIEEE_Float_1484_1908: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier1484WeightOutput, flopocoMultiplier1484WeightOutput);

    MB_D_FF_Float_1484_1908_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier1484WeightOutput, flopocoMultiplier1484WeightInput);

    MB_D_FF_Float_Multiplier9_1536_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier388_Output_492, mb_D_FFMultiplier9_1536_0Output);

    MB_D_FF_Float_1536_1971_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier9_1536_0Output, mb_D_FF1536_1971MultiplierStage1Output);

    MB_D_FF_Float_1536_1971_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1536_1971MultiplierStage1Output, mb_D_FF1536_1971MultiplierStage2Output);

    Multiplier_Float_1536: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF1536_1971MultiplierStage2Output, flopocoMultiplier1536WeightInput, Multiplier1536_Output_1971);

    MBRightSHR_Float_1536_1971: entity work.MBRightSHR(rtl)
    GENERIC MAP (160, NumberOfBits)
    PORT MAP (clk, rst, Multiplier1536Weight, mbRightSHR1536_1971Output);

    MB_D_FF_Float_1536_1971_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR1536_1971Output, Multiplier1536WeightOutput);

    InputIEEE_Float_1536_1971: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier1536WeightOutput, flopocoMultiplier1536WeightOutput);

    MB_D_FF_Float_1536_1971_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier1536WeightOutput, flopocoMultiplier1536WeightInput);

    MB_D_FF_Float_Adder8_Input1_435_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier1536_Output_1971, mb_D_FFAdder8_Input1_435_0Output);

    MB_D_FF_Float_435_1972_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder8_Input1_435_0Output, mb_D_FF435_1972AugendStage1Output);

    MB_D_FF_Float_435_1972_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF435_1972AugendStage1Output, mb_D_FF435_1972AugendStage2Output);

    Adder_Float_435: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF435_1972AugendStage2Output, mb_D_FF435_1972AddendStage2Output, Adder435_Output_1972);

    MB_D_FF_Float_Adder8_Input2_435_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier1484_Output_1908, mb_D_FFAdder8_Input2_435_0Output);

    MB_D_FF_Float_435_1972_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder8_Input2_435_0Output, mb_D_FF435_1972AddendStage1Output);

    MB_D_FF_Float_435_1972_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF435_1972AddendStage1Output, mb_D_FF435_1972AddendStage2Output);

    MB_D_FF_Float_Multiplier7_1537_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder435_Output_1972, mb_D_FFMultiplier7_1537_0Output);

    MB_D_FF_Float_1537_1973_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier7_1537_0Output, mb_D_FF1537_1973MultiplierStage1Output);

    MB_D_FF_Float_1537_1973_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1537_1973MultiplierStage1Output, mb_D_FF1537_1973MultiplierStage2Output);

    Multiplier_Float_1537: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF1537_1973MultiplierStage2Output, mb_D_FF1537_1973MultiplicandStage2Output, Multiplier1537_Output_1973);

    MBRightSHR_Float_1537_1973: entity work.MBRightSHR(rtl)
    GENERIC MAP (174, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR1537_1973Input, mbRightSHR1537_1973Output);

    MB_D_FF_Float_1537_1973_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR1537_1973Output, mb_D_FF1537_1973MultiplicandStage1Output);

    MB_D_FF_Float_1537_1973_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1537_1973MultiplicandStage1Output, mb_D_FF1537_1973MultiplicandStage2Output);

    MB_D_FF_Float_Multiplier8_1627_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier1340_Output_1723, mb_D_FFMultiplier8_1627_0Output);

    MB_D_FF_Float_1627_2092_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier8_1627_0Output, mb_D_FF1627_2092MultiplierStage1Output);

    MB_D_FF_Float_1627_2092_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1627_2092MultiplierStage1Output, mb_D_FF1627_2092MultiplierStage2Output);

    Multiplier_Float_1627: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF1627_2092MultiplierStage2Output, flopocoMultiplier1627WeightInput, Multiplier1627_Output_2092);

    MBRightSHR_Float_1627_2092: entity work.MBRightSHR(rtl)
    GENERIC MAP (167, NumberOfBits)
    PORT MAP (clk, rst, Multiplier1627Weight, mbRightSHR1627_2092Output);

    MB_D_FF_Float_1627_2092_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR1627_2092Output, Multiplier1627WeightOutput);

    InputIEEE_Float_1627_2092: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier1627WeightOutput, flopocoMultiplier1627WeightOutput);

    MB_D_FF_Float_1627_2092_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier1627WeightOutput, flopocoMultiplier1627WeightInput);

    MB_D_FF_Float_Multiplier8_1717_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier1430_Output_1842, mb_D_FFMultiplier8_1717_0Output);

    MB_D_FF_Float_1717_2211_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier8_1717_0Output, mb_D_FF1717_2211MultiplierStage1Output);

    MB_D_FF_Float_1717_2211_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1717_2211MultiplierStage1Output, mb_D_FF1717_2211MultiplierStage2Output);

    Multiplier_Float_1717: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF1717_2211MultiplierStage2Output, flopocoMultiplier1717WeightInput, Multiplier1717_Output_2211);

    MBRightSHR_Float_1717_2211: entity work.MBRightSHR(rtl)
    GENERIC MAP (167, NumberOfBits)
    PORT MAP (clk, rst, Multiplier1717Weight, mbRightSHR1717_2211Output);

    MB_D_FF_Float_1717_2211_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR1717_2211Output, Multiplier1717WeightOutput);

    InputIEEE_Float_1717_2211: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier1717WeightOutput, flopocoMultiplier1717WeightOutput);

    MB_D_FF_Float_1717_2211_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier1717WeightOutput, flopocoMultiplier1717WeightInput);

    MB_D_FF_Float_Adder7_Input1_494_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier1717_Output_2211, mb_D_FFAdder7_Input1_494_0Output);

    MB_D_FF_Float_494_2212_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder7_Input1_494_0Output, mb_D_FF494_2212AugendStage1Output);

    MB_D_FF_Float_494_2212_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF494_2212AugendStage1Output, mb_D_FF494_2212AugendStage2Output);

    Adder_Float_494: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF494_2212AugendStage2Output, mb_D_FF494_2212AddendStage2Output, Adder494_Output_2212);

    MB_D_FF_Float_Adder7_Input2_494_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier1627_Output_2092, mb_D_FFAdder7_Input2_494_0Output);

    MB_D_FF_Float_494_2212_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder7_Input2_494_0Output, mb_D_FF494_2212AddendStage1Output);

    MB_D_FF_Float_494_2212_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF494_2212AddendStage1Output, mb_D_FF494_2212AddendStage2Output);

    MB_D_FF_Float_Multiplier6_Input1_1718_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder494_Output_2212, mb_D_FFMultiplier6_Input1_1718_0Output);

    MB_D_FF_Float_1718_2213_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier6_Input1_1718_0Output, mb_D_FF1718_2213MultiplicandStage1Output);

    MB_D_FF_Float_1718_2213_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1718_2213MultiplicandStage1Output, mb_D_FF1718_2213MultiplicandStage2Output);

    Multiplier_Float_1718: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF1718_2213MultiplicandStage2Output, mb_D_FF1718_2213MultiplierStage2Output, Multiplier1718_Output_2213);

    MB_D_FF_Float_Multiplier6_Input2_1718_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier1537_Output_1973, mb_D_FFMultiplier6_Input2_1718_0Output);

    MB_D_FF_Float_1718_2213_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier6_Input2_1718_0Output, mb_D_FF1718_2213MultiplierStage1Output);

    MB_D_FF_Float_1718_2213_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1718_2213MultiplierStage1Output, mb_D_FF1718_2213MultiplierStage2Output);

    MB_D_FF_Float_Adder5_Input1_495_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier1718_Output_2213, mb_D_FFAdder5_Input1_495_0Output);

    MB_D_FF_Float_495_2214_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder5_Input1_495_0Output, mb_D_FF495_2214AugendStage1Output);

    MB_D_FF_Float_495_2214_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF495_2214AugendStage1Output, mb_D_FF495_2214AugendStage2Output);

    Adder_Float_495: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF495_2214AugendStage2Output, mb_D_FF495_2214AddendStage2Output, Adder495_Output_2214);

    MB_D_FF_Float_Adder5_Input2_495_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier1432_Output_1845, mb_D_FFAdder5_Input2_495_0Output);

    MB_D_FF_Float_495_2214_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder5_Input2_495_0Output, mb_D_FF495_2214AddendStage1Output);

    MB_D_FF_Float_495_2214_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF495_2214AddendStage1Output, mb_D_FF495_2214AddendStage2Output);

    MB_D_FF_Float_Multiplier4_1719_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder495_Output_2214, mb_D_FFMultiplier4_1719_0Output);

    MB_D_FF_Float_1719_2215_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier4_1719_0Output, mb_D_FF1719_2215MultiplierStage1Output);

    MB_D_FF_Float_1719_2215_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1719_2215MultiplierStage1Output, mb_D_FF1719_2215MultiplierStage2Output);

    Multiplier_Float_1719: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF1719_2215MultiplierStage2Output, mb_D_FF1719_2215MultiplicandStage2Output, Multiplier1719_Output_2215);

    MBRightSHR_Float_1719_2215: entity work.MBRightSHR(rtl)
    GENERIC MAP (231, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR1719_2215Input, mbRightSHR1719_2215Output);

    MB_D_FF_Float_1719_2215_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR1719_2215Output, mb_D_FF1719_2215MultiplicandStage1Output);

    MB_D_FF_Float_1719_2215_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1719_2215MultiplicandStage1Output, mb_D_FF1719_2215MultiplicandStage2Output);

    MB_D_FF_Float_Multiplier9_1771_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier623_Output_799, mb_D_FFMultiplier9_1771_0Output);

    MB_D_FF_Float_1771_2278_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier9_1771_0Output, mb_D_FF1771_2278MultiplierStage1Output);

    MB_D_FF_Float_1771_2278_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1771_2278MultiplierStage1Output, mb_D_FF1771_2278MultiplierStage2Output);

    Multiplier_Float_1771: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF1771_2278MultiplierStage2Output, flopocoMultiplier1771WeightInput, Multiplier1771_Output_2278);

    MBRightSHR_Float_1771_2278: entity work.MBRightSHR(rtl)
    GENERIC MAP (160, NumberOfBits)
    PORT MAP (clk, rst, Multiplier1771Weight, mbRightSHR1771_2278Output);

    MB_D_FF_Float_1771_2278_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR1771_2278Output, Multiplier1771WeightOutput);

    InputIEEE_Float_1771_2278: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier1771WeightOutput, flopocoMultiplier1771WeightOutput);

    MB_D_FF_Float_1771_2278_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier1771WeightOutput, flopocoMultiplier1771WeightInput);

    MB_D_FF_Float_Multiplier9_1823_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier675_Output_862, mb_D_FFMultiplier9_1823_0Output);

    MB_D_FF_Float_1823_2341_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier9_1823_0Output, mb_D_FF1823_2341MultiplierStage1Output);

    MB_D_FF_Float_1823_2341_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1823_2341MultiplierStage1Output, mb_D_FF1823_2341MultiplierStage2Output);

    Multiplier_Float_1823: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF1823_2341MultiplierStage2Output, flopocoMultiplier1823WeightInput, Multiplier1823_Output_2341);

    MBRightSHR_Float_1823_2341: entity work.MBRightSHR(rtl)
    GENERIC MAP (160, NumberOfBits)
    PORT MAP (clk, rst, Multiplier1823Weight, mbRightSHR1823_2341Output);

    MB_D_FF_Float_1823_2341_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR1823_2341Output, Multiplier1823WeightOutput);

    InputIEEE_Float_1823_2341: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier1823WeightOutput, flopocoMultiplier1823WeightOutput);

    MB_D_FF_Float_1823_2341_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier1823WeightOutput, flopocoMultiplier1823WeightInput);

    MB_D_FF_Float_Adder8_Input1_518_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier1823_Output_2341, mb_D_FFAdder8_Input1_518_0Output);

    MB_D_FF_Float_518_2342_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder8_Input1_518_0Output, mb_D_FF518_2342AugendStage1Output);

    MB_D_FF_Float_518_2342_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF518_2342AugendStage1Output, mb_D_FF518_2342AugendStage2Output);

    Adder_Float_518: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF518_2342AugendStage2Output, mb_D_FF518_2342AddendStage2Output, Adder518_Output_2342);

    MB_D_FF_Float_Adder8_Input2_518_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier1771_Output_2278, mb_D_FFAdder8_Input2_518_0Output);

    MB_D_FF_Float_518_2342_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder8_Input2_518_0Output, mb_D_FF518_2342AddendStage1Output);

    MB_D_FF_Float_518_2342_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF518_2342AddendStage1Output, mb_D_FF518_2342AddendStage2Output);

    MB_D_FF_Float_Multiplier7_1824_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder518_Output_2342, mb_D_FFMultiplier7_1824_0Output);

    MB_D_FF_Float_1824_2343_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier7_1824_0Output, mb_D_FF1824_2343MultiplierStage1Output);

    MB_D_FF_Float_1824_2343_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1824_2343MultiplierStage1Output, mb_D_FF1824_2343MultiplierStage2Output);

    Multiplier_Float_1824: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF1824_2343MultiplierStage2Output, mb_D_FF1824_2343MultiplicandStage2Output, Multiplier1824_Output_2343);

    MBRightSHR_Float_1824_2343: entity work.MBRightSHR(rtl)
    GENERIC MAP (174, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR1824_2343Input, mbRightSHR1824_2343Output);

    MB_D_FF_Float_1824_2343_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR1824_2343Output, mb_D_FF1824_2343MultiplicandStage1Output);

    MB_D_FF_Float_1824_2343_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1824_2343MultiplicandStage1Output, mb_D_FF1824_2343MultiplicandStage2Output);

    MB_D_FF_Float_Multiplier11_Input1_1868_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder367_Output_1662, mb_D_FFMultiplier11_Input1_1868_0Output);

    MB_D_FF_Float_1868_2401_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier11_Input1_1868_0Output, mb_D_FF1868_2401MultiplicandStage1Output);

    MB_D_FF_Float_1868_2401_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1868_2401MultiplicandStage1Output, mb_D_FF1868_2401MultiplicandStage2Output);

    Multiplier_Float_1868: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF1868_2401MultiplicandStage2Output, mb_D_FF1868_2401MultiplierStage2Output, Multiplier1868_Output_2401);

    MB_D_FF_Float_Multiplier11_Input2_1868_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier710_Output_909, mb_D_FFMultiplier11_Input2_1868_0Output);

    MB_D_FF_Float_1868_2401_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier11_Input2_1868_0Output, mb_D_FF1868_2401MultiplierStage1Output);

    MB_D_FF_Float_1868_2401_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1868_2401MultiplierStage1Output, mb_D_FF1868_2401MultiplierStage2Output);

    MB_D_FF_Float_Multiplier11_Input1_1912_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder381_Output_1720, mb_D_FFMultiplier11_Input1_1912_0Output);

    MB_D_FF_Float_1912_2459_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier11_Input1_1912_0Output, mb_D_FF1912_2459MultiplicandStage1Output);

    MB_D_FF_Float_1912_2459_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1912_2459MultiplicandStage1Output, mb_D_FF1912_2459MultiplicandStage2Output);

    Multiplier_Float_1912: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF1912_2459MultiplicandStage2Output, mb_D_FF1912_2459MultiplierStage2Output, Multiplier1912_Output_2459);

    MB_D_FF_Float_Multiplier11_Input2_1912_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier754_Output_967, mb_D_FFMultiplier11_Input2_1912_0Output);

    MB_D_FF_Float_1912_2459_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier11_Input2_1912_0Output, mb_D_FF1912_2459MultiplierStage1Output);

    MB_D_FF_Float_1912_2459_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1912_2459MultiplierStage1Output, mb_D_FF1912_2459MultiplierStage2Output);

    MB_D_FF_Float_Adder10_Input1_547_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier1912_Output_2459, mb_D_FFAdder10_Input1_547_0Output);

    MB_D_FF_Float_547_2460_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder10_Input1_547_0Output, mb_D_FF547_2460AugendStage1Output);

    MB_D_FF_Float_547_2460_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF547_2460AugendStage1Output, mb_D_FF547_2460AugendStage2Output);

    Adder_Float_547: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF547_2460AugendStage2Output, mb_D_FF547_2460AddendStage2Output, Adder547_Output_2460);

    MB_D_FF_Float_Adder10_Input2_547_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier1868_Output_2401, mb_D_FFAdder10_Input2_547_0Output);

    MB_D_FF_Float_547_2460_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder10_Input2_547_0Output, mb_D_FF547_2460AddendStage1Output);

    MB_D_FF_Float_547_2460_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF547_2460AddendStage1Output, mb_D_FF547_2460AddendStage2Output);

    MB_D_FF_Float_Multiplier9_1913_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder547_Output_2460, mb_D_FFMultiplier9_1913_0Output);

    MB_D_FF_Float_1913_2461_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier9_1913_0Output, mb_D_FF1913_2461MultiplierStage1Output);

    MB_D_FF_Float_1913_2461_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1913_2461MultiplierStage1Output, mb_D_FF1913_2461MultiplierStage2Output);

    Multiplier_Float_1913: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF1913_2461MultiplierStage2Output, mb_D_FF1913_2461MultiplicandStage2Output, Multiplier1913_Output_2461);

    MBRightSHR_Float_1913_2461: entity work.MBRightSHR(rtl)
    GENERIC MAP (160, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR1913_2461Input, mbRightSHR1913_2461Output);

    MB_D_FF_Float_1913_2461_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR1913_2461Output, mb_D_FF1913_2461MultiplicandStage1Output);

    MB_D_FF_Float_1913_2461_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1913_2461MultiplicandStage1Output, mb_D_FF1913_2461MultiplicandStage2Output);

    MB_D_FF_Float_Multiplier8_1914_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier1913_Output_2461, mb_D_FFMultiplier8_1914_0Output);

    MB_D_FF_Float_1914_2462_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier8_1914_0Output, mb_D_FF1914_2462MultiplierStage1Output);

    MB_D_FF_Float_1914_2462_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1914_2462MultiplierStage1Output, mb_D_FF1914_2462MultiplierStage2Output);

    Multiplier_Float_1914: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF1914_2462MultiplierStage2Output, flopocoMultiplier1914WeightInput, Multiplier1914_Output_2462);

    MBRightSHR_Float_1914_2462: entity work.MBRightSHR(rtl)
    GENERIC MAP (167, NumberOfBits)
    PORT MAP (clk, rst, Multiplier1914Weight, mbRightSHR1914_2462Output);

    MB_D_FF_Float_1914_2462_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR1914_2462Output, Multiplier1914WeightOutput);

    InputIEEE_Float_1914_2462: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier1914WeightOutput, flopocoMultiplier1914WeightOutput);

    MB_D_FF_Float_1914_2462_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier1914WeightOutput, flopocoMultiplier1914WeightInput);

    MB_D_FF_Float_Multiplier11_Input1_1958_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder396_Output_1781, mb_D_FFMultiplier11_Input1_1958_0Output);

    MB_D_FF_Float_1958_2520_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier11_Input1_1958_0Output, mb_D_FF1958_2520MultiplicandStage1Output);

    MB_D_FF_Float_1958_2520_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1958_2520MultiplicandStage1Output, mb_D_FF1958_2520MultiplicandStage2Output);

    Multiplier_Float_1958: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF1958_2520MultiplicandStage2Output, mb_D_FF1958_2520MultiplierStage2Output, Multiplier1958_Output_2520);

    MB_D_FF_Float_Multiplier11_Input2_1958_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier800_Output_1028, mb_D_FFMultiplier11_Input2_1958_0Output);

    MB_D_FF_Float_1958_2520_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier11_Input2_1958_0Output, mb_D_FF1958_2520MultiplierStage1Output);

    MB_D_FF_Float_1958_2520_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1958_2520MultiplierStage1Output, mb_D_FF1958_2520MultiplierStage2Output);

    MB_D_FF_Float_Multiplier11_Input1_2002_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder410_Output_1839, mb_D_FFMultiplier11_Input1_2002_0Output);

    MB_D_FF_Float_2002_2578_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier11_Input1_2002_0Output, mb_D_FF2002_2578MultiplicandStage1Output);

    MB_D_FF_Float_2002_2578_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF2002_2578MultiplicandStage1Output, mb_D_FF2002_2578MultiplicandStage2Output);

    Multiplier_Float_2002: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF2002_2578MultiplicandStage2Output, mb_D_FF2002_2578MultiplierStage2Output, Multiplier2002_Output_2578);

    MB_D_FF_Float_Multiplier11_Input2_2002_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier844_Output_1086, mb_D_FFMultiplier11_Input2_2002_0Output);

    MB_D_FF_Float_2002_2578_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier11_Input2_2002_0Output, mb_D_FF2002_2578MultiplierStage1Output);

    MB_D_FF_Float_2002_2578_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF2002_2578MultiplierStage1Output, mb_D_FF2002_2578MultiplierStage2Output);

    MB_D_FF_Float_Adder10_Input1_576_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier2002_Output_2578, mb_D_FFAdder10_Input1_576_0Output);

    MB_D_FF_Float_576_2579_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder10_Input1_576_0Output, mb_D_FF576_2579AugendStage1Output);

    MB_D_FF_Float_576_2579_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF576_2579AugendStage1Output, mb_D_FF576_2579AugendStage2Output);

    Adder_Float_576: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF576_2579AugendStage2Output, mb_D_FF576_2579AddendStage2Output, Adder576_Output_2579);

    MB_D_FF_Float_Adder10_Input2_576_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier1958_Output_2520, mb_D_FFAdder10_Input2_576_0Output);

    MB_D_FF_Float_576_2579_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder10_Input2_576_0Output, mb_D_FF576_2579AddendStage1Output);

    MB_D_FF_Float_576_2579_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF576_2579AddendStage1Output, mb_D_FF576_2579AddendStage2Output);

    MB_D_FF_Float_Multiplier9_2003_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder576_Output_2579, mb_D_FFMultiplier9_2003_0Output);

    MB_D_FF_Float_2003_2580_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier9_2003_0Output, mb_D_FF2003_2580MultiplierStage1Output);

    MB_D_FF_Float_2003_2580_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF2003_2580MultiplierStage1Output, mb_D_FF2003_2580MultiplierStage2Output);

    Multiplier_Float_2003: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF2003_2580MultiplierStage2Output, mb_D_FF2003_2580MultiplicandStage2Output, Multiplier2003_Output_2580);

    MBRightSHR_Float_2003_2580: entity work.MBRightSHR(rtl)
    GENERIC MAP (160, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR2003_2580Input, mbRightSHR2003_2580Output);

    MB_D_FF_Float_2003_2580_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR2003_2580Output, mb_D_FF2003_2580MultiplicandStage1Output);

    MB_D_FF_Float_2003_2580_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF2003_2580MultiplicandStage1Output, mb_D_FF2003_2580MultiplicandStage2Output);

    MB_D_FF_Float_Multiplier8_2004_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier2003_Output_2580, mb_D_FFMultiplier8_2004_0Output);

    MB_D_FF_Float_2004_2581_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier8_2004_0Output, mb_D_FF2004_2581MultiplierStage1Output);

    MB_D_FF_Float_2004_2581_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF2004_2581MultiplierStage1Output, mb_D_FF2004_2581MultiplierStage2Output);

    Multiplier_Float_2004: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF2004_2581MultiplierStage2Output, flopocoMultiplier2004WeightInput, Multiplier2004_Output_2581);

    MBRightSHR_Float_2004_2581: entity work.MBRightSHR(rtl)
    GENERIC MAP (167, NumberOfBits)
    PORT MAP (clk, rst, Multiplier2004Weight, mbRightSHR2004_2581Output);

    MB_D_FF_Float_2004_2581_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR2004_2581Output, Multiplier2004WeightOutput);

    InputIEEE_Float_2004_2581: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier2004WeightOutput, flopocoMultiplier2004WeightOutput);

    MB_D_FF_Float_2004_2581_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier2004WeightOutput, flopocoMultiplier2004WeightInput);

    MB_D_FF_Float_Adder7_Input1_577_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier2004_Output_2581, mb_D_FFAdder7_Input1_577_0Output);

    MB_D_FF_Float_577_2582_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder7_Input1_577_0Output, mb_D_FF577_2582AugendStage1Output);

    MB_D_FF_Float_577_2582_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF577_2582AugendStage1Output, mb_D_FF577_2582AugendStage2Output);

    Adder_Float_577: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF577_2582AugendStage2Output, mb_D_FF577_2582AddendStage2Output, Adder577_Output_2582);

    MB_D_FF_Float_Adder7_Input2_577_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier1914_Output_2462, mb_D_FFAdder7_Input2_577_0Output);

    MB_D_FF_Float_577_2582_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder7_Input2_577_0Output, mb_D_FF577_2582AddendStage1Output);

    MB_D_FF_Float_577_2582_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF577_2582AddendStage1Output, mb_D_FF577_2582AddendStage2Output);

    MB_D_FF_Float_Multiplier6_Input1_2005_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder577_Output_2582, mb_D_FFMultiplier6_Input1_2005_0Output);

    MB_D_FF_Float_2005_2583_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier6_Input1_2005_0Output, mb_D_FF2005_2583MultiplicandStage1Output);

    MB_D_FF_Float_2005_2583_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF2005_2583MultiplicandStage1Output, mb_D_FF2005_2583MultiplicandStage2Output);

    Multiplier_Float_2005: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF2005_2583MultiplicandStage2Output, mb_D_FF2005_2583MultiplierStage2Output, Multiplier2005_Output_2583);

    MB_D_FF_Float_Multiplier6_Input2_2005_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier1824_Output_2343, mb_D_FFMultiplier6_Input2_2005_0Output);

    MB_D_FF_Float_2005_2583_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier6_Input2_2005_0Output, mb_D_FF2005_2583MultiplierStage1Output);

    MB_D_FF_Float_2005_2583_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF2005_2583MultiplierStage1Output, mb_D_FF2005_2583MultiplierStage2Output);

    MB_D_FF_Float_Multiplier9_2057_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier909_Output_1167, mb_D_FFMultiplier9_2057_0Output);

    MB_D_FF_Float_2057_2646_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier9_2057_0Output, mb_D_FF2057_2646MultiplierStage1Output);

    MB_D_FF_Float_2057_2646_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF2057_2646MultiplierStage1Output, mb_D_FF2057_2646MultiplierStage2Output);

    Multiplier_Float_2057: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF2057_2646MultiplierStage2Output, flopocoMultiplier2057WeightInput, Multiplier2057_Output_2646);

    MBRightSHR_Float_2057_2646: entity work.MBRightSHR(rtl)
    GENERIC MAP (160, NumberOfBits)
    PORT MAP (clk, rst, Multiplier2057Weight, mbRightSHR2057_2646Output);

    MB_D_FF_Float_2057_2646_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR2057_2646Output, Multiplier2057WeightOutput);

    InputIEEE_Float_2057_2646: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier2057WeightOutput, flopocoMultiplier2057WeightOutput);

    MB_D_FF_Float_2057_2646_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier2057WeightOutput, flopocoMultiplier2057WeightInput);

    MB_D_FF_Float_Multiplier9_2109_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier961_Output_1230, mb_D_FFMultiplier9_2109_0Output);

    MB_D_FF_Float_2109_2709_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier9_2109_0Output, mb_D_FF2109_2709MultiplierStage1Output);

    MB_D_FF_Float_2109_2709_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF2109_2709MultiplierStage1Output, mb_D_FF2109_2709MultiplierStage2Output);

    Multiplier_Float_2109: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF2109_2709MultiplierStage2Output, flopocoMultiplier2109WeightInput, Multiplier2109_Output_2709);

    MBRightSHR_Float_2109_2709: entity work.MBRightSHR(rtl)
    GENERIC MAP (160, NumberOfBits)
    PORT MAP (clk, rst, Multiplier2109Weight, mbRightSHR2109_2709Output);

    MB_D_FF_Float_2109_2709_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR2109_2709Output, Multiplier2109WeightOutput);

    InputIEEE_Float_2109_2709: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier2109WeightOutput, flopocoMultiplier2109WeightOutput);

    MB_D_FF_Float_2109_2709_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier2109WeightOutput, flopocoMultiplier2109WeightInput);

    MB_D_FF_Float_Adder8_Input1_600_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier2109_Output_2709, mb_D_FFAdder8_Input1_600_0Output);

    MB_D_FF_Float_600_2710_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder8_Input1_600_0Output, mb_D_FF600_2710AugendStage1Output);

    MB_D_FF_Float_600_2710_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF600_2710AugendStage1Output, mb_D_FF600_2710AugendStage2Output);

    Adder_Float_600: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF600_2710AugendStage2Output, mb_D_FF600_2710AddendStage2Output, Adder600_Output_2710);

    MB_D_FF_Float_Adder8_Input2_600_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier2057_Output_2646, mb_D_FFAdder8_Input2_600_0Output);

    MB_D_FF_Float_600_2710_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder8_Input2_600_0Output, mb_D_FF600_2710AddendStage1Output);

    MB_D_FF_Float_600_2710_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF600_2710AddendStage1Output, mb_D_FF600_2710AddendStage2Output);

    MB_D_FF_Float_Multiplier7_2110_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder600_Output_2710, mb_D_FFMultiplier7_2110_0Output);

    MB_D_FF_Float_2110_2711_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier7_2110_0Output, mb_D_FF2110_2711MultiplierStage1Output);

    MB_D_FF_Float_2110_2711_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF2110_2711MultiplierStage1Output, mb_D_FF2110_2711MultiplierStage2Output);

    Multiplier_Float_2110: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF2110_2711MultiplierStage2Output, mb_D_FF2110_2711MultiplicandStage2Output, Multiplier2110_Output_2711);

    MBRightSHR_Float_2110_2711: entity work.MBRightSHR(rtl)
    GENERIC MAP (174, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR2110_2711Input, mbRightSHR2110_2711Output);

    MB_D_FF_Float_2110_2711_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR2110_2711Output, mb_D_FF2110_2711MultiplicandStage1Output);

    MB_D_FF_Float_2110_2711_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF2110_2711MultiplicandStage1Output, mb_D_FF2110_2711MultiplicandStage2Output);

    MB_D_FF_Float_Multiplier8_2200_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier1913_Output_2461, mb_D_FFMultiplier8_2200_0Output);

    MB_D_FF_Float_2200_2830_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier8_2200_0Output, mb_D_FF2200_2830MultiplierStage1Output);

    MB_D_FF_Float_2200_2830_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF2200_2830MultiplierStage1Output, mb_D_FF2200_2830MultiplierStage2Output);

    Multiplier_Float_2200: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF2200_2830MultiplierStage2Output, flopocoMultiplier2200WeightInput, Multiplier2200_Output_2830);

    MBRightSHR_Float_2200_2830: entity work.MBRightSHR(rtl)
    GENERIC MAP (167, NumberOfBits)
    PORT MAP (clk, rst, Multiplier2200Weight, mbRightSHR2200_2830Output);

    MB_D_FF_Float_2200_2830_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR2200_2830Output, Multiplier2200WeightOutput);

    InputIEEE_Float_2200_2830: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier2200WeightOutput, flopocoMultiplier2200WeightOutput);

    MB_D_FF_Float_2200_2830_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier2200WeightOutput, flopocoMultiplier2200WeightInput);

    MB_D_FF_Float_Multiplier8_2290_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier2003_Output_2580, mb_D_FFMultiplier8_2290_0Output);

    MB_D_FF_Float_2290_2949_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier8_2290_0Output, mb_D_FF2290_2949MultiplierStage1Output);

    MB_D_FF_Float_2290_2949_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF2290_2949MultiplierStage1Output, mb_D_FF2290_2949MultiplierStage2Output);

    Multiplier_Float_2290: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF2290_2949MultiplierStage2Output, flopocoMultiplier2290WeightInput, Multiplier2290_Output_2949);

    MBRightSHR_Float_2290_2949: entity work.MBRightSHR(rtl)
    GENERIC MAP (167, NumberOfBits)
    PORT MAP (clk, rst, Multiplier2290Weight, mbRightSHR2290_2949Output);

    MB_D_FF_Float_2290_2949_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR2290_2949Output, Multiplier2290WeightOutput);

    InputIEEE_Float_2290_2949: entity work.InputIEEE_7_14_to_7_14(arch)
        PORT MAP (clk, Multiplier2290WeightOutput, flopocoMultiplier2290WeightOutput);

    MB_D_FF_Float_2290_2949_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier2290WeightOutput, flopocoMultiplier2290WeightInput);

    MB_D_FF_Float_Adder7_Input1_659_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier2290_Output_2949, mb_D_FFAdder7_Input1_659_0Output);

    MB_D_FF_Float_659_2950_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder7_Input1_659_0Output, mb_D_FF659_2950AugendStage1Output);

    MB_D_FF_Float_659_2950_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF659_2950AugendStage1Output, mb_D_FF659_2950AugendStage2Output);

    Adder_Float_659: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF659_2950AugendStage2Output, mb_D_FF659_2950AddendStage2Output, Adder659_Output_2950);

    MB_D_FF_Float_Adder7_Input2_659_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier2200_Output_2830, mb_D_FFAdder7_Input2_659_0Output);

    MB_D_FF_Float_659_2950_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder7_Input2_659_0Output, mb_D_FF659_2950AddendStage1Output);

    MB_D_FF_Float_659_2950_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF659_2950AddendStage1Output, mb_D_FF659_2950AddendStage2Output);

    MB_D_FF_Float_Multiplier6_Input1_2291_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder659_Output_2950, mb_D_FFMultiplier6_Input1_2291_0Output);

    MB_D_FF_Float_2291_2951_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier6_Input1_2291_0Output, mb_D_FF2291_2951MultiplicandStage1Output);

    MB_D_FF_Float_2291_2951_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF2291_2951MultiplicandStage1Output, mb_D_FF2291_2951MultiplicandStage2Output);

    Multiplier_Float_2291: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF2291_2951MultiplicandStage2Output, mb_D_FF2291_2951MultiplierStage2Output, Multiplier2291_Output_2951);

    MB_D_FF_Float_Multiplier6_Input2_2291_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier2110_Output_2711, mb_D_FFMultiplier6_Input2_2291_0Output);

    MB_D_FF_Float_2291_2951_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier6_Input2_2291_0Output, mb_D_FF2291_2951MultiplierStage1Output);

    MB_D_FF_Float_2291_2951_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF2291_2951MultiplierStage1Output, mb_D_FF2291_2951MultiplierStage2Output);

    MB_D_FF_Float_Adder5_Input1_660_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier2291_Output_2951, mb_D_FFAdder5_Input1_660_0Output);

    MB_D_FF_Float_660_2952_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder5_Input1_660_0Output, mb_D_FF660_2952AugendStage1Output);

    MB_D_FF_Float_660_2952_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF660_2952AugendStage1Output, mb_D_FF660_2952AugendStage2Output);

    Adder_Float_660: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF660_2952AugendStage2Output, mb_D_FF660_2952AddendStage2Output, Adder660_Output_2952);

    MB_D_FF_Float_Adder5_Input2_660_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier2005_Output_2583, mb_D_FFAdder5_Input2_660_0Output);

    MB_D_FF_Float_660_2952_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder5_Input2_660_0Output, mb_D_FF660_2952AddendStage1Output);

    MB_D_FF_Float_660_2952_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF660_2952AddendStage1Output, mb_D_FF660_2952AddendStage2Output);

    MB_D_FF_Float_Multiplier4_2292_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder660_Output_2952, mb_D_FFMultiplier4_2292_0Output);

    MB_D_FF_Float_2292_2953_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier4_2292_0Output, mb_D_FF2292_2953MultiplierStage1Output);

    MB_D_FF_Float_2292_2953_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF2292_2953MultiplierStage1Output, mb_D_FF2292_2953MultiplierStage2Output);

    Multiplier_Float_2292: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF2292_2953MultiplierStage2Output, mb_D_FF2292_2953MultiplicandStage2Output, Multiplier2292_Output_2953);

    MBRightSHR_Float_2292_2953: entity work.MBRightSHR(rtl)
    GENERIC MAP (231, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR2292_2953Input, mbRightSHR2292_2953Output);

    MB_D_FF_Float_2292_2953_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR2292_2953Output, mb_D_FF2292_2953MultiplicandStage1Output);

    MB_D_FF_Float_2292_2953_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF2292_2953MultiplicandStage1Output, mb_D_FF2292_2953MultiplicandStage2Output);

    MB_D_FF_Float_Adder3_Input1_661_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier2292_Output_2953, mb_D_FFAdder3_Input1_661_0Output);

    MB_D_FF_Float_661_2954_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder3_Input1_661_0Output, mb_D_FF661_2954AugendStage1Output);

    MB_D_FF_Float_661_2954_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF661_2954AugendStage1Output, mb_D_FF661_2954AugendStage2Output);

    Adder_Float_661: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF661_2954AugendStage2Output, mb_D_FF661_2954AddendStage2Output, Adder661_Output_2954);

    MB_D_FF_Float_Adder3_Input2_661_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier1719_Output_2215, mb_D_FFAdder3_Input2_661_0Output);

    MB_D_FF_Float_661_2954_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder3_Input2_661_0Output, mb_D_FF661_2954AddendStage1Output);

    MB_D_FF_Float_661_2954_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF661_2954AddendStage1Output, mb_D_FF661_2954AddendStage2Output);

    MB_D_FF_Float_Multiplier2_2293_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder661_Output_2954, mb_D_FFMultiplier2_2293_0Output);

    MB_D_FF_Float_2293_2955_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier2_2293_0Output, mb_D_FF2293_2955MultiplierStage1Output);

    MB_D_FF_Float_2293_2955_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF2293_2955MultiplierStage1Output, mb_D_FF2293_2955MultiplierStage2Output);

    Multiplier_Float_2293: entity work.FPMult_7_14_7_14_7_14_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF2293_2955MultiplierStage2Output, mb_D_FF2293_2955MultiplicandStage2Output, Multiplier2293_Output_2955);

    MBRightSHR_Float_2293_2955: entity work.MBRightSHR(rtl)
    GENERIC MAP (263, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR2293_2955Input, mbRightSHR2293_2955Output);

    MB_D_FF_Float_2293_2955_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR2293_2955Output, mb_D_FF2293_2955MultiplicandStage1Output);

    MB_D_FF_Float_2293_2955_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF2293_2955MultiplicandStage1Output, mb_D_FF2293_2955MultiplicandStage2Output);

    MB_D_FF_Float_Adder1_Input1_662_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier2293_Output_2955, mb_D_FFAdder1_Input1_662_0Output);

    MB_D_FF_Float_662_2956_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder1_Input1_662_0Output, mb_D_FF662_2956AugendStage1Output);

    MB_D_FF_Float_662_2956_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF662_2956AugendStage1Output, mb_D_FF662_2956AugendStage2Output);

    Adder_Float_662: entity work.FPAdd_7_14_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF662_2956AugendStage2Output, mb_D_FF662_2956AddendStage2Output, Adder662_Output_2956);

    MB_D_FF_Float_Adder1_Input2_662_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier1146_Output_1477, mb_D_FFAdder1_Input2_662_0Output);

    MB_D_FF_Float_662_2956_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder1_Input2_662_0Output, mb_D_FF662_2956AddendStage1Output);

    MB_D_FF_Float_662_2956_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF662_2956AddendStage1Output, mb_D_FF662_2956AddendStage2Output);

    MB_D_FF_Float_Adder1_Output_662_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder662_Output_2956, mb_D_FFAdder1_Output_662_0Output);

    vout <= mb_D_FFAdder1_Output_662_0Output;
 
END ARCHITECTURE;

LIBRARY ieee; 
LIBRARY ieee_proposed; 
USE ieee.std_logic_1164.all; 
USE ieee.std_logic_arith.all; 
USE ieee.std_logic_unsigned.all; 
USE ieee.std_logic_textio.all; 
 
LIBRARY std; 
USE std.textio.all; 
USE ieee_proposed.fixed_pkg.all; 
USE ieee_proposed.fixed_float_types.all; 
USE ieee_proposed.float_pkg.all; 
ENTITY PCSystem_32 IS
    GENERIC (MantissaBits :INTEGER := 25 ; ExponentBits :INTEGER := 7 ; NumberOfBits :INTEGER := 32 ; FlopocoBits :INTEGER := 2);
    PORT (
    clk:IN std_logic;
    rst:IN std_logic;
    enable:IN std_logic;
    v0a:IN std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
    v0b:IN std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
    v1a:IN std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
    v1b:IN std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
    v2a:IN std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
    v2b:IN std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
    v3a:IN std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
    v3b:IN std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
    v4a:IN std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
    v4b:IN std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
    v5a:IN std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
    v5b:IN std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
    v6a:IN std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
    v6b:IN std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
    v7a:IN std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
    v7b:IN std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
    v8a:IN std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
    v8b:IN std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
    v9a:IN std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
    v9b:IN std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
    v10a:IN std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
    v10b:IN std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
    v11a:IN std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
    v11b:IN std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
    v12a:IN std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
    v12b:IN std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
    v13a:IN std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
    v13b:IN std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
    v14a:IN std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
    v14b:IN std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
    v15a:IN std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
    v15b:IN std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
    v16a:IN std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
    v16b:IN std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
    vout:OUT std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0)
);
END PCSystem_32;

ARCHITECTURE rtl of PCSystem_32 IS

        SIGNAL mb_D_FFMultiplier2_102_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier102_Output_136 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier102WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier102WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier102WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF102_136MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF102_136MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR102_136Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier2_53_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier53_Output_71 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier53WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier53WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier53WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF53_71MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF53_71MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR53_71Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier3_101_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier101_Output_135 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF101_135MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF101_135MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF101_135MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF101_135MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR101_135Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR101_135Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier3_Input1_52_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier52_Output_70 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF52_70MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF52_70MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF52_70MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF52_70MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier3_Input2_52_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier4_Input1_100_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier100_Output_134 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF100_134MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF100_134MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF100_134MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF100_134MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier4_Input2_100_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder4_Input1_17_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder17_Output_69 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF17_69AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF17_69AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF17_69AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF17_69AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder4_Input2_17_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier4_Input1_49_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier49_Output_66 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF49_66MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF49_66MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF49_66MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF49_66MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier4_Input2_49_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder5_Input1_33_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder33_Output_133 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF33_133AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF33_133AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF33_133AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF33_133AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder5_Input2_33_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier5_Input1_97_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier97_Output_130 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF97_130MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF97_130MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF97_130MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF97_130MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier5_Input2_97_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier51_Output_68 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier51WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier51WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier51WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF51_68MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF51_68MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR51_Input1_68Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR51_Input2_68Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR51_Input2_68Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier50_Output_67 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier50WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier50WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier50WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF50_67MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF50_67MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR50_Input1_67Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR50_Input2_67Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR50_Input2_67Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder5_Input1_16_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder16_Output_65 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF16_65AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF16_65AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF16_65AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF16_65AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder5_Input2_16_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier5_Input1_46_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier46_Output_62 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF46_62MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF46_62MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF46_62MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF46_62MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier5_Input2_46_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier99_Output_132 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier99WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier99WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier99WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF99_132MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF99_132MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR99_Input1_132Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR99_Input2_132Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR99_Input2_132Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier98_Output_131 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier98WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier98WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier98WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF98_131MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF98_131MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR98_Input1_131Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR98_Input2_131Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR98_Input2_131Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder6_Input1_32_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder32_Output_129 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF32_129AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF32_129AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF32_129AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF32_129AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder6_Input2_32_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier6_Input1_94_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier94_Output_126 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF94_126MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF94_126MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF94_126MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF94_126MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier6_Input2_94_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier48_Output_64 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier48WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier48WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier48WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF48_64MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF48_64MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR48_Input1_64Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR48_Input2_64Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR48_Input2_64Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier47_Output_63 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier47WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier47WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier47WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF47_63MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF47_63MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR47_Input1_63Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR47_Input2_63Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR47_Input2_63Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder6_Input1_15_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder15_Output_61 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF15_61AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF15_61AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF15_61AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF15_61AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder6_Input2_15_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier6_Input1_43_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier43_Output_58 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF43_58MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF43_58MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF43_58MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF43_58MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier6_Input2_43_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier96_Output_128 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier96WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier96WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier96WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF96_128MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF96_128MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR96_Input1_128Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR96_Input2_128Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR96_Input2_128Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier95_Output_127 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier95WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier95WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier95WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF95_127MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF95_127MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR95_Input1_127Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR95_Input2_127Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR95_Input2_127Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder7_Input1_31_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder31_Output_125 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF31_125AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF31_125AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF31_125AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF31_125AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder7_Input2_31_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier7_Input1_91_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier91_Output_122 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF91_122MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF91_122MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF91_122MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF91_122MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier7_Input2_91_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier45_Output_60 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier45WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier45WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier45WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF45_60MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF45_60MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR45_Input1_60Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR45_Input2_60Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR45_Input2_60Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier44_Output_59 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier44WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier44WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier44WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF44_59MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF44_59MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR44_Input1_59Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR44_Input2_59Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR44_Input2_59Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder7_Input1_14_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder14_Output_57 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF14_57AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF14_57AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF14_57AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF14_57AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder7_Input2_14_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier7_Input1_40_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier40_Output_54 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF40_54MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF40_54MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF40_54MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF40_54MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier7_Input2_40_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier93_Output_124 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier93WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier93WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier93WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF93_124MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF93_124MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR93_Input1_124Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR93_Input2_124Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR93_Input2_124Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier92_Output_123 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier92WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier92WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier92WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF92_123MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF92_123MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR92_Input1_123Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR92_Input2_123Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR92_Input2_123Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder8_Input1_30_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder30_Output_121 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF30_121AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF30_121AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF30_121AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF30_121AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder8_Input2_30_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier8_Input1_88_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier88_Output_118 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF88_118MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF88_118MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF88_118MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF88_118MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier8_Input2_88_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier42_Output_56 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier42WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier42WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier42WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF42_56MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF42_56MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR42_Input1_56Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR42_Input2_56Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR42_Input2_56Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier41_Output_55 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier41WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier41WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier41WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF41_55MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF41_55MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR41_Input1_55Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR41_Input2_55Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR41_Input2_55Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder8_Input1_13_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder13_Output_53 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF13_53AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF13_53AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF13_53AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF13_53AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder8_Input2_13_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier8_Input1_37_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier37_Output_50 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF37_50MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF37_50MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF37_50MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF37_50MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier8_Input2_37_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier90_Output_120 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier90WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier90WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier90WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF90_120MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF90_120MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR90_Input1_120Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR90_Input2_120Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR90_Input2_120Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier89_Output_119 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier89WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier89WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier89WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF89_119MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF89_119MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR89_Input1_119Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR89_Input2_119Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR89_Input2_119Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder9_Input1_29_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder29_Output_117 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF29_117AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF29_117AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF29_117AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF29_117AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder9_Input2_29_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier9_Input1_85_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier85_Output_114 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF85_114MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF85_114MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF85_114MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF85_114MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier9_Input2_85_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier39_Output_52 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier39WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier39WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier39WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF39_52MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF39_52MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR39_Input1_52Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR39_Input2_52Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR39_Input2_52Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier38_Output_51 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier38WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier38WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier38WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF38_51MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF38_51MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR38_Input1_51Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR38_Input2_51Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR38_Input2_51Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder9_Input1_12_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder12_Output_49 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF12_49AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF12_49AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF12_49AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF12_49AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder9_Input2_12_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier9_Input1_34_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier34_Output_46 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF34_46MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF34_46MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF34_46MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF34_46MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier9_Input2_34_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier87_Output_116 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier87WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier87WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier87WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF87_116MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF87_116MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR87_Input1_116Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR87_Input2_116Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR87_Input2_116Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier86_Output_115 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier86WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier86WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier86WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF86_115MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF86_115MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR86_Input1_115Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR86_Input2_115Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR86_Input2_115Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder10_Input1_28_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder28_Output_113 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF28_113AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF28_113AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF28_113AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF28_113AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder10_Input2_28_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier10_Input1_82_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier82_Output_110 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF82_110MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF82_110MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF82_110MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF82_110MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier10_Input2_82_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier36_Output_48 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier36WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier36WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier36WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF36_48MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF36_48MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR36_Input1_48Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR36_Input2_48Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR36_Input2_48Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier35_Output_47 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier35WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier35WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier35WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF35_47MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF35_47MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR35_Input1_47Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR35_Input2_47Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR35_Input2_47Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder10_Input1_11_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder11_Output_45 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF11_45AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF11_45AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF11_45AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF11_45AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder10_Input2_11_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier10_Input1_31_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier31_Output_42 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF31_42MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF31_42MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF31_42MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF31_42MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier10_Input2_31_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier84_Output_112 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier84WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier84WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier84WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF84_112MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF84_112MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR84_Input1_112Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR84_Input2_112Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR84_Input2_112Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier83_Output_111 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier83WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier83WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier83WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF83_111MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF83_111MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR83_Input1_111Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR83_Input2_111Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR83_Input2_111Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder11_Input1_27_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder27_Output_109 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF27_109AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF27_109AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF27_109AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF27_109AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder11_Input2_27_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier11_Input1_79_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier79_Output_106 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF79_106MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF79_106MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF79_106MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF79_106MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier11_Input2_79_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier33_Output_44 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier33WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier33WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier33WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF33_44MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF33_44MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR33_Input1_44Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR33_Input2_44Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR33_Input2_44Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier32_Output_43 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier32WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier32WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier32WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF32_43MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF32_43MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR32_Input1_43Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR32_Input2_43Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR32_Input2_43Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder11_Input1_10_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder10_Output_41 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF10_41AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF10_41AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF10_41AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF10_41AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder11_Input2_10_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier11_Input1_28_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier28_Output_38 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF28_38MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF28_38MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF28_38MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF28_38MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier11_Input2_28_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier81_Output_108 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier81WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier81WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier81WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF81_108MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF81_108MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR81_Input1_108Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR81_Input2_108Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR81_Input2_108Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier80_Output_107 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier80WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier80WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier80WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF80_107MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF80_107MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR80_Input1_107Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR80_Input2_107Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR80_Input2_107Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder12_Input1_26_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder26_Output_105 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF26_105AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF26_105AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF26_105AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF26_105AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder12_Input2_26_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier12_Input1_76_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier76_Output_102 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF76_102MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF76_102MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF76_102MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF76_102MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier12_Input2_76_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier30_Output_40 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier30WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier30WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier30WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF30_40MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF30_40MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR30_Input1_40Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR30_Input2_40Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR30_Input2_40Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier29_Output_39 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier29WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier29WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier29WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF29_39MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF29_39MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR29_Input1_39Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR29_Input2_39Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR29_Input2_39Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder12_Input1_9_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder9_Output_37 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF9_37AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF9_37AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF9_37AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF9_37AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder12_Input2_9_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier12_Input1_25_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier25_Output_34 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF25_34MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF25_34MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF25_34MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF25_34MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier12_Input2_25_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier78_Output_104 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier78WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier78WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier78WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF78_104MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF78_104MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR78_Input1_104Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR78_Input2_104Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR78_Input2_104Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier77_Output_103 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier77WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier77WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier77WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF77_103MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF77_103MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR77_Input1_103Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR77_Input2_103Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR77_Input2_103Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder13_Input1_25_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder25_Output_101 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF25_101AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF25_101AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF25_101AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF25_101AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder13_Input2_25_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier13_Input1_73_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier73_Output_98 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF73_98MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF73_98MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF73_98MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF73_98MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier13_Input2_73_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier27_Output_36 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier27WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier27WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier27WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF27_36MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF27_36MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR27_Input1_36Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR27_Input2_36Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR27_Input2_36Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier26_Output_35 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier26WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier26WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier26WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF26_35MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF26_35MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR26_Input1_35Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR26_Input2_35Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR26_Input2_35Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder13_Input1_8_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder8_Output_33 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF8_33AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF8_33AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF8_33AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF8_33AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder13_Input2_8_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier13_Input1_22_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier22_Output_30 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF22_30MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF22_30MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF22_30MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF22_30MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier13_Input2_22_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier75_Output_100 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier75WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier75WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier75WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF75_100MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF75_100MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR75_Input1_100Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR75_Input2_100Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR75_Input2_100Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier74_Output_99 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier74WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier74WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier74WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF74_99MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF74_99MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR74_Input1_99Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR74_Input2_99Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR74_Input2_99Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder14_Input1_24_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder24_Output_97 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF24_97AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF24_97AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF24_97AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF24_97AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder14_Input2_24_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier14_Input1_70_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier70_Output_94 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF70_94MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF70_94MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF70_94MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF70_94MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier14_Input2_70_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier24_Output_32 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier24WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier24WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier24WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF24_32MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF24_32MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR24_Input1_32Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR24_Input2_32Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR24_Input2_32Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier23_Output_31 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier23WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier23WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier23WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF23_31MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF23_31MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR23_Input1_31Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR23_Input2_31Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR23_Input2_31Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder14_Input1_7_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder7_Output_29 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF7_29AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF7_29AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF7_29AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF7_29AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder14_Input2_7_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier14_Input1_19_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier19_Output_26 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF19_26MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF19_26MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF19_26MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF19_26MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier14_Input2_19_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier72_Output_96 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier72WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier72WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier72WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF72_96MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF72_96MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR72_Input1_96Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR72_Input2_96Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR72_Input2_96Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier71_Output_95 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier71WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier71WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier71WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF71_95MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF71_95MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR71_Input1_95Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR71_Input2_95Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR71_Input2_95Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder15_Input1_23_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder23_Output_93 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF23_93AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF23_93AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF23_93AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF23_93AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder15_Input2_23_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier15_Input1_67_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier67_Output_90 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF67_90MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF67_90MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF67_90MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF67_90MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier15_Input2_67_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier21_Output_28 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier21WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier21WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier21WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF21_28MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF21_28MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR21_Input1_28Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR21_Input2_28Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR21_Input2_28Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier20_Output_27 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier20WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier20WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier20WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF20_27MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF20_27MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR20_Input1_27Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR20_Input2_27Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR20_Input2_27Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder15_Input1_6_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder6_Output_25 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF6_25AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF6_25AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF6_25AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF6_25AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder15_Input2_6_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier15_Input1_16_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier16_Output_22 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF16_22MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF16_22MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF16_22MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF16_22MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier15_Input2_16_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier69_Output_92 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier69WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier69WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier69WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF69_92MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF69_92MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR69_Input1_92Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR69_Input2_92Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR69_Input2_92Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier68_Output_91 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier68WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier68WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier68WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF68_91MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF68_91MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR68_Input1_91Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR68_Input2_91Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR68_Input2_91Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder16_Input1_22_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder22_Output_89 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF22_89AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF22_89AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF22_89AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF22_89AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder16_Input2_22_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier16_Input1_64_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier64_Output_86 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF64_86MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF64_86MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF64_86MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF64_86MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier16_Input2_64_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier18_Output_24 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier18WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier18WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier18WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF18_24MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF18_24MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR18_Input1_24Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR18_Input2_24Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR18_Input2_24Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier17_Output_23 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier17WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier17WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier17WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF17_23MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF17_23MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR17_Input1_23Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR17_Input2_23Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR17_Input2_23Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder16_Input1_5_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder5_Output_21 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF5_21AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF5_21AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF5_21AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF5_21AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder16_Input2_5_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier16_Input1_7_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier7_Output_10 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF7_10MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF7_10MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF7_10MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF7_10MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier16_Input2_7_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier66_Output_88 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier66WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier66WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier66WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF66_88MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF66_88MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR66_Input1_88Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR66_Input2_88Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR66_Input2_88Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier65_Output_87 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier65WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier65WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier65WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF65_87MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF65_87MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR65_Input1_87Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR65_Input2_87Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR65_Input2_87Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder17_Input1_21_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder21_Output_85 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF21_85AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF21_85AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF21_85AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF21_85AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder17_Input2_21_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier17_Input1_61_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier61_Output_82 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF61_82MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF61_82MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF61_82MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF61_82MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier17_Input2_61_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier17_15_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier15_Output_20 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier15WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier15WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier15WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF15_20MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF15_20MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR15_20Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier17_11_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier11_Output_15 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier11WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier11WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier11WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF11_15MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF11_15MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR11_15Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFAdder17_Input1_2_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder2_Output_9 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF2_9AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF2_9AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF2_9AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF2_9AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder17_Input2_2_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier17_Input1_4_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier4_Output_6 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF4_6MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF4_6MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF4_6MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF4_6MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier17_Input2_4_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier63_Output_84 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier63WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier63WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier63WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF63_84MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF63_84MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR63_Input1_84Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR63_Input2_84Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR63_Input2_84Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier62_Output_83 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier62WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier62WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier62WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF62_83MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF62_83MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR62_Input1_83Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR62_Input2_83Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR62_Input2_83Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder18_Input1_20_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder20_Output_81 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF20_81AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF20_81AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF20_81AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF20_81AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder18_Input2_20_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier18_Input1_58_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier58_Output_78 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF58_78MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF58_78MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF58_78MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF58_78MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier18_Input2_58_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier18_14_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier14_Output_19 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF14_19MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF14_19MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF14_19MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF14_19MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR14_19Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR14_19Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier18_10_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier10_Output_14 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF10_14MultiplicandStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF10_14MultiplicandStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF10_14MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF10_14MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR10_14Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR10_14Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier6_Output_8 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier6WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier6WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier6WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF6_8MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF6_8MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR6_Input1_8Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR6_Input2_8Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR6_Input2_8Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier5_Output_7 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier5WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier5WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier5WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF5_7MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF5_7MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR5_Input1_7Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR5_Input2_7Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR5_Input2_7Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder18_Input1_1_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder1_Output_5 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1_5AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1_5AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1_5AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1_5AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder18_Input2_1_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder18_Input1_0_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder0_Output_2 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF0_2AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF0_2AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF0_2AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF0_2AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder18_Input2_0_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier60_Output_80 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier60WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier60WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier60WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF60_80MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF60_80MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR60_Input1_80Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR60_Input2_80Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR60_Input2_80Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier59_Output_79 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier59WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier59WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier59WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF59_79MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF59_79MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR59_Input1_79Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR59_Input2_79Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR59_Input2_79Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder19_Input1_19_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder19_Output_77 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF19_77AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF19_77AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF19_77AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF19_77AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder19_Input2_19_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder19_Input1_18_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder18_Output_74 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF18_74AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF18_74AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF18_74AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF18_74AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder19_Input2_18_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder19_Input1_4_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder4_Output_18 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF4_18AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF4_18AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF4_18AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF4_18AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder19_Input2_4_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder19_Input1_3_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder3_Output_13 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF3_13AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF3_13AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF3_13AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF3_13AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder19_Input2_3_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier3_Output_4 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier3WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier3WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier3WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF3_4MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF3_4MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR3_Input1_4Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR3_Input2_4Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR3_Input2_4Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier2_Output_3 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier2WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier2WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier2WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF2_3MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF2_3MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR2_Input1_3Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR2_Input2_3Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR2_Input2_3Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1_Output_1 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier1WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier1WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier1WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1_1MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF1_1MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1_Input1_1Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR1_Input2_1Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR1_Input2_1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier0_Output_0 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier0WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier0WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier0WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF0_0MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF0_0MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR0_Input1_0Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mbRightSHR0_Input2_0Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR0_Input2_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier57_Output_76 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier57WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier57WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier57WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF57_76MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF57_76MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR57_76Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier20_57_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier20_57_0Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier56_Output_75 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier56WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier56WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier56WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF56_75MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF56_75MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR56_75Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier20_56_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier20_56_0Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier55_Output_73 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier55WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier55WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier55WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF55_73MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF55_73MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR55_73Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier20_55_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier20_55_0Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier54_Output_72 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier54WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier54WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier54WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF54_72MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF54_72MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR54_72Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier20_54_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier20_54_0Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier13_Output_17 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier13WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier13WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier13WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF13_17MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF13_17MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR13_17Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier20_13_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier20_13_0Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier12_Output_16 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier12WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier12WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier12WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF12_16MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF12_16MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR12_16Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier20_12_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier20_12_0Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier9_Output_12 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier9WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier9WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier9WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF9_12MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF9_12MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR9_12Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier20_9_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier20_9_0Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier8_Output_11 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL flopocoMultiplier8WeightOutput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier8WeightOutput :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL flopocoMultiplier8WeightInput :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF8_11MultiplierStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF8_11MultiplierStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mbRightSHR8_11Output :std_logic_vector(NumberOfBits-1 DOWNTO 0);

        SIGNAL mb_D_FFMultiplier20_8_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFMultiplier20_8_0Input :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder1_Input1_34_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Adder34_Output_137 :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF34_137AugendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF34_137AugendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF34_137AddendStage1Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FF34_137AddendStage2Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder1_Input2_34_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL mb_D_FFAdder1_Output_34_0Output :std_logic_vector(FlopocoBits+(MantissaBits-1)+(ExponentBits) DOWNTO 0);
        SIGNAL Multiplier0Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.013664569414715357,exponentBits,mantissaBits-1));
        SIGNAL Multiplier1Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.9863354305852846,exponentBits,mantissaBits-1));
        SIGNAL Multiplier2Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.0031062391443788602,exponentBits,mantissaBits-1));
        SIGNAL Multiplier3Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.9968937608556211,exponentBits,mantissaBits-1));
        SIGNAL Multiplier5Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.0849999639647431,exponentBits,mantissaBits-1));
        SIGNAL Multiplier6Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.9150000360352569,exponentBits,mantissaBits-1));
        SIGNAL Multiplier8Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.4438857309430112,exponentBits,mantissaBits-1));
        SIGNAL Multiplier9Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.5561142690569888,exponentBits,mantissaBits-1));
        SIGNAL Multiplier11Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.19779031804717737,exponentBits,mantissaBits-1));
        SIGNAL Multiplier12Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.1167201214636732,exponentBits,mantissaBits-1));
        SIGNAL Multiplier13Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.8832798785363268,exponentBits,mantissaBits-1));
        SIGNAL Multiplier15Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.8022096819528226,exponentBits,mantissaBits-1));
        SIGNAL Multiplier17Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.15583807196961508,exponentBits,mantissaBits-1));
        SIGNAL Multiplier18Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.8441619280303849,exponentBits,mantissaBits-1));
        SIGNAL Multiplier20Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.082491910084827,exponentBits,mantissaBits-1));
        SIGNAL Multiplier21Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.917508089915173,exponentBits,mantissaBits-1));
        SIGNAL Multiplier23Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.08289550496205488,exponentBits,mantissaBits-1));
        SIGNAL Multiplier24Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.9171044950379451,exponentBits,mantissaBits-1));
        SIGNAL Multiplier26Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.25200175852053647,exponentBits,mantissaBits-1));
        SIGNAL Multiplier27Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.7479982414794635,exponentBits,mantissaBits-1));
        SIGNAL Multiplier29Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.15867765021296837,exponentBits,mantissaBits-1));
        SIGNAL Multiplier30Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.8413223497870317,exponentBits,mantissaBits-1));
        SIGNAL Multiplier32Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.7638321333592787,exponentBits,mantissaBits-1));
        SIGNAL Multiplier33Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.2361678666407213,exponentBits,mantissaBits-1));
        SIGNAL Multiplier35Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.36282458757648484,exponentBits,mantissaBits-1));
        SIGNAL Multiplier36Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.6371754124235152,exponentBits,mantissaBits-1));
        SIGNAL Multiplier38Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.05344749302717779,exponentBits,mantissaBits-1));
        SIGNAL Multiplier39Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.9465525069728222,exponentBits,mantissaBits-1));
        SIGNAL Multiplier41Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.2661492003776495,exponentBits,mantissaBits-1));
        SIGNAL Multiplier42Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.7338507996223504,exponentBits,mantissaBits-1));
        SIGNAL Multiplier44Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.19119586603532895,exponentBits,mantissaBits-1));
        SIGNAL Multiplier45Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.808804133964671,exponentBits,mantissaBits-1));
        SIGNAL Multiplier47Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.2404344410571303,exponentBits,mantissaBits-1));
        SIGNAL Multiplier48Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.7595655589428697,exponentBits,mantissaBits-1));
        SIGNAL Multiplier50Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.0007639474461813438,exponentBits,mantissaBits-1));
        SIGNAL Multiplier51Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.9992360525538186,exponentBits,mantissaBits-1));
        SIGNAL Multiplier53Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.47628086748179016,exponentBits,mantissaBits-1));
        SIGNAL Multiplier54Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.03718220130691538,exponentBits,mantissaBits-1));
        SIGNAL Multiplier55Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.9628177986930846,exponentBits,mantissaBits-1));
        SIGNAL Multiplier56Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.006187202191737726,exponentBits,mantissaBits-1));
        SIGNAL Multiplier57Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.9938127978082623,exponentBits,mantissaBits-1));
        SIGNAL Multiplier59Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.04552574833030746,exponentBits,mantissaBits-1));
        SIGNAL Multiplier60Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.9544742516696926,exponentBits,mantissaBits-1));
        SIGNAL Multiplier62Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.8093371697482517,exponentBits,mantissaBits-1));
        SIGNAL Multiplier63Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.19066283025174835,exponentBits,mantissaBits-1));
        SIGNAL Multiplier65Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.01829288275120762,exponentBits,mantissaBits-1));
        SIGNAL Multiplier66Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.9817071172487923,exponentBits,mantissaBits-1));
        SIGNAL Multiplier68Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.21115138327226968,exponentBits,mantissaBits-1));
        SIGNAL Multiplier69Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.7888486167277303,exponentBits,mantissaBits-1));
        SIGNAL Multiplier71Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.16135227071631283,exponentBits,mantissaBits-1));
        SIGNAL Multiplier72Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.8386477292836871,exponentBits,mantissaBits-1));
        SIGNAL Multiplier74Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.1291709542317448,exponentBits,mantissaBits-1));
        SIGNAL Multiplier75Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.8708290457682553,exponentBits,mantissaBits-1));
        SIGNAL Multiplier77Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.05495074488933167,exponentBits,mantissaBits-1));
        SIGNAL Multiplier78Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.9450492551106683,exponentBits,mantissaBits-1));
        SIGNAL Multiplier80Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.05257811015055088,exponentBits,mantissaBits-1));
        SIGNAL Multiplier81Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.9474218898494491,exponentBits,mantissaBits-1));
        SIGNAL Multiplier83Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.17826220890983333,exponentBits,mantissaBits-1));
        SIGNAL Multiplier84Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.8217377910901666,exponentBits,mantissaBits-1));
        SIGNAL Multiplier86Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.19620771696171668,exponentBits,mantissaBits-1));
        SIGNAL Multiplier87Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.8037922830382833,exponentBits,mantissaBits-1));
        SIGNAL Multiplier89Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.060266233212953796,exponentBits,mantissaBits-1));
        SIGNAL Multiplier90Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.9397337667870462,exponentBits,mantissaBits-1));
        SIGNAL Multiplier92Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.19243902918602898,exponentBits,mantissaBits-1));
        SIGNAL Multiplier93Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.807560970813971,exponentBits,mantissaBits-1));
        SIGNAL Multiplier95Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.1636790257778244,exponentBits,mantissaBits-1));
        SIGNAL Multiplier96Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.8363209742221756,exponentBits,mantissaBits-1));
        SIGNAL Multiplier98Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.36697842999744384,exponentBits,mantissaBits-1));
        SIGNAL Multiplier99Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.6330215700025561,exponentBits,mantissaBits-1));
        SIGNAL Multiplier102Weight :std_logic_vector(NumberOfBits-1 DOWNTO 0):= to_slv(to_float(0.5237191325182098,exponentBits,mantissaBits-1));
        
BEGIN
    PROCESS (clk,rst) IS
    BEGIN 
        IF rst = '1' THEN
    mbRightSHR101_135Input <= (others=>'0');
mbRightSHR51_Input2_68Input <= (others=>'0');
            mbRightSHR50_Input2_67Input <= (others=>'0');
mbRightSHR99_Input2_132Input <= (others=>'0');
            mbRightSHR98_Input2_131Input <= (others=>'0');
            mbRightSHR48_Input2_64Input <= (others=>'0');
            mbRightSHR47_Input2_63Input <= (others=>'0');
mbRightSHR96_Input2_128Input <= (others=>'0');
            mbRightSHR95_Input2_127Input <= (others=>'0');
            mbRightSHR45_Input2_60Input <= (others=>'0');
            mbRightSHR44_Input2_59Input <= (others=>'0');
mbRightSHR93_Input2_124Input <= (others=>'0');
            mbRightSHR92_Input2_123Input <= (others=>'0');
            mbRightSHR42_Input2_56Input <= (others=>'0');
            mbRightSHR41_Input2_55Input <= (others=>'0');
mbRightSHR90_Input2_120Input <= (others=>'0');
            mbRightSHR89_Input2_119Input <= (others=>'0');
            mbRightSHR39_Input2_52Input <= (others=>'0');
            mbRightSHR38_Input2_51Input <= (others=>'0');
mbRightSHR87_Input2_116Input <= (others=>'0');
            mbRightSHR86_Input2_115Input <= (others=>'0');
            mbRightSHR36_Input2_48Input <= (others=>'0');
            mbRightSHR35_Input2_47Input <= (others=>'0');
mbRightSHR84_Input2_112Input <= (others=>'0');
            mbRightSHR83_Input2_111Input <= (others=>'0');
            mbRightSHR33_Input2_44Input <= (others=>'0');
            mbRightSHR32_Input2_43Input <= (others=>'0');
mbRightSHR81_Input2_108Input <= (others=>'0');
            mbRightSHR80_Input2_107Input <= (others=>'0');
            mbRightSHR30_Input2_40Input <= (others=>'0');
            mbRightSHR29_Input2_39Input <= (others=>'0');
mbRightSHR78_Input2_104Input <= (others=>'0');
            mbRightSHR77_Input2_103Input <= (others=>'0');
            mbRightSHR27_Input2_36Input <= (others=>'0');
            mbRightSHR26_Input2_35Input <= (others=>'0');
mbRightSHR75_Input2_100Input <= (others=>'0');
            mbRightSHR74_Input2_99Input <= (others=>'0');
            mbRightSHR24_Input2_32Input <= (others=>'0');
            mbRightSHR23_Input2_31Input <= (others=>'0');
mbRightSHR72_Input2_96Input <= (others=>'0');
            mbRightSHR71_Input2_95Input <= (others=>'0');
            mbRightSHR21_Input2_28Input <= (others=>'0');
            mbRightSHR20_Input2_27Input <= (others=>'0');
mbRightSHR69_Input2_92Input <= (others=>'0');
            mbRightSHR68_Input2_91Input <= (others=>'0');
            mbRightSHR18_Input2_24Input <= (others=>'0');
            mbRightSHR17_Input2_23Input <= (others=>'0');
mbRightSHR66_Input2_88Input <= (others=>'0');
            mbRightSHR65_Input2_87Input <= (others=>'0');
mbRightSHR63_Input2_84Input <= (others=>'0');
            mbRightSHR62_Input2_83Input <= (others=>'0');
            mbRightSHR14_19Input <= (others=>'0');
            mbRightSHR10_14Input <= (others=>'0');
            mbRightSHR6_Input2_8Input <= (others=>'0');
            mbRightSHR5_Input2_7Input <= (others=>'0');
mbRightSHR60_Input2_80Input <= (others=>'0');
            mbRightSHR59_Input2_79Input <= (others=>'0');
            mbRightSHR3_Input2_4Input <= (others=>'0');
            mbRightSHR2_Input2_3Input <= (others=>'0');
            mbRightSHR1_Input2_1Input <= (others=>'0');
            mbRightSHR0_Input2_0Input <= (others=>'0');
mb_D_FFMultiplier20_57_0Input <= (others=>'0');
            mb_D_FFMultiplier20_56_0Input <= (others=>'0');
            mb_D_FFMultiplier20_55_0Input <= (others=>'0');
            mb_D_FFMultiplier20_54_0Input <= (others=>'0');
            mb_D_FFMultiplier20_13_0Input <= (others=>'0');
            mb_D_FFMultiplier20_12_0Input <= (others=>'0');
            mb_D_FFMultiplier20_9_0Input <= (others=>'0');
            mb_D_FFMultiplier20_8_0Input <= (others=>'0');
        ELSIF rising_edge(clk) and rst = '0' and enable = '1' THEN
            mbRightSHR101_135Input <= v0b;
mbRightSHR51_Input2_68Input <= v0a;
            mbRightSHR50_Input2_67Input <= v0b;
mbRightSHR99_Input2_132Input <= v1a;
            mbRightSHR98_Input2_131Input <= v1b;
            mbRightSHR48_Input2_64Input <= v1a;
            mbRightSHR47_Input2_63Input <= v1b;
mbRightSHR96_Input2_128Input <= v2a;
            mbRightSHR95_Input2_127Input <= v2b;
            mbRightSHR45_Input2_60Input <= v2a;
            mbRightSHR44_Input2_59Input <= v2b;
mbRightSHR93_Input2_124Input <= v3a;
            mbRightSHR92_Input2_123Input <= v3b;
            mbRightSHR42_Input2_56Input <= v3a;
            mbRightSHR41_Input2_55Input <= v3b;
mbRightSHR90_Input2_120Input <= v4a;
            mbRightSHR89_Input2_119Input <= v4b;
            mbRightSHR39_Input2_52Input <= v4a;
            mbRightSHR38_Input2_51Input <= v4b;
mbRightSHR87_Input2_116Input <= v5a;
            mbRightSHR86_Input2_115Input <= v5b;
            mbRightSHR36_Input2_48Input <= v5a;
            mbRightSHR35_Input2_47Input <= v5b;
mbRightSHR84_Input2_112Input <= v6a;
            mbRightSHR83_Input2_111Input <= v6b;
            mbRightSHR33_Input2_44Input <= v6b;
            mbRightSHR32_Input2_43Input <= v6a;
mbRightSHR81_Input2_108Input <= v7a;
            mbRightSHR80_Input2_107Input <= v7b;
            mbRightSHR30_Input2_40Input <= v7a;
            mbRightSHR29_Input2_39Input <= v7b;
mbRightSHR78_Input2_104Input <= v8a;
            mbRightSHR77_Input2_103Input <= v8b;
            mbRightSHR27_Input2_36Input <= v8a;
            mbRightSHR26_Input2_35Input <= v8b;
mbRightSHR75_Input2_100Input <= v9a;
            mbRightSHR74_Input2_99Input <= v9b;
            mbRightSHR24_Input2_32Input <= v9a;
            mbRightSHR23_Input2_31Input <= v9b;
mbRightSHR72_Input2_96Input <= v10a;
            mbRightSHR71_Input2_95Input <= v10b;
            mbRightSHR21_Input2_28Input <= v10a;
            mbRightSHR20_Input2_27Input <= v10b;
mbRightSHR69_Input2_92Input <= v11a;
            mbRightSHR68_Input2_91Input <= v11b;
            mbRightSHR18_Input2_24Input <= v11a;
            mbRightSHR17_Input2_23Input <= v11b;
mbRightSHR66_Input2_88Input <= v12a;
            mbRightSHR65_Input2_87Input <= v12b;
mbRightSHR63_Input2_84Input <= v13b;
            mbRightSHR62_Input2_83Input <= v13a;
            mbRightSHR14_19Input <= v13a;
            mbRightSHR10_14Input <= v13b;
            mbRightSHR6_Input2_8Input <= v14a;
            mbRightSHR5_Input2_7Input <= v14b;
mbRightSHR60_Input2_80Input <= v14a;
            mbRightSHR59_Input2_79Input <= v14b;
            mbRightSHR3_Input2_4Input <= v15a;
            mbRightSHR2_Input2_3Input <= v15b;
            mbRightSHR1_Input2_1Input <= v16a;
            mbRightSHR0_Input2_0Input <= v16b;
mb_D_FFMultiplier20_57_0Input <= v15a;
            mb_D_FFMultiplier20_56_0Input <= v15b;
            mb_D_FFMultiplier20_55_0Input <= v16a;
            mb_D_FFMultiplier20_54_0Input <= v16b;
            mb_D_FFMultiplier20_13_0Input <= v12a;
            mb_D_FFMultiplier20_12_0Input <= v12b;
            mb_D_FFMultiplier20_9_0Input <= v12a;
            mb_D_FFMultiplier20_8_0Input <= v12b;
        END IF;

    END PROCESS;

    MBRightSHR_Float_0_Input10: entity work.MBRightSHR(rtl)
    GENERIC MAP (16, NumberOfBits)
    PORT MAP (clk, rst, Multiplier0Weight, mbRightSHR0_Input1_0Output);

    MB_D_FF_Float_0_0_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR0_Input1_0Output, Multiplier0WeightOutput);

    InputIEEE_Float_0_0: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier0WeightOutput, flopocoMultiplier0WeightOutput);

    MB_D_FF_Float_0_0_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier0WeightOutput, flopocoMultiplier0WeightInput);

    Multiplier_Float_0: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier0WeightInput, mb_D_FF0_0MultiplierStage2Output, Multiplier0_Output_0);

    MBRightSHR_Float_0_Input2_0: entity work.MBRightSHR(rtl)
    GENERIC MAP (16, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR0_Input2_0Input, mbRightSHR0_Input2_0Output);

    MB_D_FF_Float_0_0_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR0_Input2_0Output, mb_D_FF0_0MultiplierStage1Output);

    MB_D_FF_Float_0_0_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF0_0MultiplierStage1Output, mb_D_FF0_0MultiplierStage2Output);

    MBRightSHR_Float_1_Input11: entity work.MBRightSHR(rtl)
    GENERIC MAP (16, NumberOfBits)
    PORT MAP (clk, rst, Multiplier1Weight, mbRightSHR1_Input1_1Output);

    MB_D_FF_Float_1_1_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR1_Input1_1Output, Multiplier1WeightOutput);

    InputIEEE_Float_1_1: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier1WeightOutput, flopocoMultiplier1WeightOutput);

    MB_D_FF_Float_1_1_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier1WeightOutput, flopocoMultiplier1WeightInput);

    Multiplier_Float_1: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier1WeightInput, mb_D_FF1_1MultiplierStage2Output, Multiplier1_Output_1);

    MBRightSHR_Float_1_Input2_1: entity work.MBRightSHR(rtl)
    GENERIC MAP (16, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR1_Input2_1Input, mbRightSHR1_Input2_1Output);

    MB_D_FF_Float_1_1_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR1_Input2_1Output, mb_D_FF1_1MultiplierStage1Output);

    MB_D_FF_Float_1_1_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1_1MultiplierStage1Output, mb_D_FF1_1MultiplierStage2Output);

    MB_D_FF_Float_Adder18_Input1_0_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier1_Output_1, mb_D_FFAdder18_Input1_0_0Output);

    MB_D_FF_Float_0_2_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder18_Input1_0_0Output, mb_D_FF0_2AugendStage1Output);

    MB_D_FF_Float_0_2_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF0_2AugendStage1Output, mb_D_FF0_2AugendStage2Output);

    Adder_Float_0: entity work.FPAdd_7_24_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF0_2AugendStage2Output, mb_D_FF0_2AddendStage2Output, Adder0_Output_2);

    MB_D_FF_Float_Adder18_Input2_0_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier0_Output_0, mb_D_FFAdder18_Input2_0_0Output);

    MB_D_FF_Float_0_2_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder18_Input2_0_0Output, mb_D_FF0_2AddendStage1Output);

    MB_D_FF_Float_0_2_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF0_2AddendStage1Output, mb_D_FF0_2AddendStage2Output);

    MBRightSHR_Float_2_Input13: entity work.MBRightSHR(rtl)
    GENERIC MAP (16, NumberOfBits)
    PORT MAP (clk, rst, Multiplier2Weight, mbRightSHR2_Input1_3Output);

    MB_D_FF_Float_2_3_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR2_Input1_3Output, Multiplier2WeightOutput);

    InputIEEE_Float_2_3: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier2WeightOutput, flopocoMultiplier2WeightOutput);

    MB_D_FF_Float_2_3_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier2WeightOutput, flopocoMultiplier2WeightInput);

    Multiplier_Float_2: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier2WeightInput, mb_D_FF2_3MultiplierStage2Output, Multiplier2_Output_3);

    MBRightSHR_Float_2_Input2_3: entity work.MBRightSHR(rtl)
    GENERIC MAP (16, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR2_Input2_3Input, mbRightSHR2_Input2_3Output);

    MB_D_FF_Float_2_3_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR2_Input2_3Output, mb_D_FF2_3MultiplierStage1Output);

    MB_D_FF_Float_2_3_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF2_3MultiplierStage1Output, mb_D_FF2_3MultiplierStage2Output);

    MBRightSHR_Float_3_Input14: entity work.MBRightSHR(rtl)
    GENERIC MAP (16, NumberOfBits)
    PORT MAP (clk, rst, Multiplier3Weight, mbRightSHR3_Input1_4Output);

    MB_D_FF_Float_3_4_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR3_Input1_4Output, Multiplier3WeightOutput);

    InputIEEE_Float_3_4: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier3WeightOutput, flopocoMultiplier3WeightOutput);

    MB_D_FF_Float_3_4_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier3WeightOutput, flopocoMultiplier3WeightInput);

    Multiplier_Float_3: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier3WeightInput, mb_D_FF3_4MultiplierStage2Output, Multiplier3_Output_4);

    MBRightSHR_Float_3_Input2_4: entity work.MBRightSHR(rtl)
    GENERIC MAP (16, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR3_Input2_4Input, mbRightSHR3_Input2_4Output);

    MB_D_FF_Float_3_4_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR3_Input2_4Output, mb_D_FF3_4MultiplierStage1Output);

    MB_D_FF_Float_3_4_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF3_4MultiplierStage1Output, mb_D_FF3_4MultiplierStage2Output);

    MB_D_FF_Float_Adder18_Input1_1_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier3_Output_4, mb_D_FFAdder18_Input1_1_0Output);

    MB_D_FF_Float_1_5_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder18_Input1_1_0Output, mb_D_FF1_5AugendStage1Output);

    MB_D_FF_Float_1_5_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1_5AugendStage1Output, mb_D_FF1_5AugendStage2Output);

    Adder_Float_1: entity work.FPAdd_7_24_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF1_5AugendStage2Output, mb_D_FF1_5AddendStage2Output, Adder1_Output_5);

    MB_D_FF_Float_Adder18_Input2_1_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier2_Output_3, mb_D_FFAdder18_Input2_1_0Output);

    MB_D_FF_Float_1_5_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder18_Input2_1_0Output, mb_D_FF1_5AddendStage1Output);

    MB_D_FF_Float_1_5_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF1_5AddendStage1Output, mb_D_FF1_5AddendStage2Output);

    MB_D_FF_Float_Multiplier17_Input1_4_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder1_Output_5, mb_D_FFMultiplier17_Input1_4_0Output);

    MB_D_FF_Float_4_6_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier17_Input1_4_0Output, mb_D_FF4_6MultiplicandStage1Output);

    MB_D_FF_Float_4_6_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF4_6MultiplicandStage1Output, mb_D_FF4_6MultiplicandStage2Output);

    Multiplier_Float_4: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF4_6MultiplicandStage2Output, mb_D_FF4_6MultiplierStage2Output, Multiplier4_Output_6);

    MB_D_FF_Float_Multiplier17_Input2_4_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder0_Output_2, mb_D_FFMultiplier17_Input2_4_0Output);

    MB_D_FF_Float_4_6_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier17_Input2_4_0Output, mb_D_FF4_6MultiplierStage1Output);

    MB_D_FF_Float_4_6_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF4_6MultiplierStage1Output, mb_D_FF4_6MultiplierStage2Output);

    MBRightSHR_Float_5_Input17: entity work.MBRightSHR(rtl)
    GENERIC MAP (43, NumberOfBits)
    PORT MAP (clk, rst, Multiplier5Weight, mbRightSHR5_Input1_7Output);

    MB_D_FF_Float_5_7_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR5_Input1_7Output, Multiplier5WeightOutput);

    InputIEEE_Float_5_7: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier5WeightOutput, flopocoMultiplier5WeightOutput);

    MB_D_FF_Float_5_7_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier5WeightOutput, flopocoMultiplier5WeightInput);

    Multiplier_Float_5: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier5WeightInput, mb_D_FF5_7MultiplierStage2Output, Multiplier5_Output_7);

    MBRightSHR_Float_5_Input2_7: entity work.MBRightSHR(rtl)
    GENERIC MAP (43, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR5_Input2_7Input, mbRightSHR5_Input2_7Output);

    MB_D_FF_Float_5_7_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR5_Input2_7Output, mb_D_FF5_7MultiplierStage1Output);

    MB_D_FF_Float_5_7_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF5_7MultiplierStage1Output, mb_D_FF5_7MultiplierStage2Output);

    MBRightSHR_Float_6_Input18: entity work.MBRightSHR(rtl)
    GENERIC MAP (43, NumberOfBits)
    PORT MAP (clk, rst, Multiplier6Weight, mbRightSHR6_Input1_8Output);

    MB_D_FF_Float_6_8_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR6_Input1_8Output, Multiplier6WeightOutput);

    InputIEEE_Float_6_8: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier6WeightOutput, flopocoMultiplier6WeightOutput);

    MB_D_FF_Float_6_8_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier6WeightOutput, flopocoMultiplier6WeightInput);

    Multiplier_Float_6: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier6WeightInput, mb_D_FF6_8MultiplierStage2Output, Multiplier6_Output_8);

    MBRightSHR_Float_6_Input2_8: entity work.MBRightSHR(rtl)
    GENERIC MAP (43, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR6_Input2_8Input, mbRightSHR6_Input2_8Output);

    MB_D_FF_Float_6_8_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR6_Input2_8Output, mb_D_FF6_8MultiplierStage1Output);

    MB_D_FF_Float_6_8_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF6_8MultiplierStage1Output, mb_D_FF6_8MultiplierStage2Output);

    MB_D_FF_Float_Adder17_Input1_2_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier6_Output_8, mb_D_FFAdder17_Input1_2_0Output);

    MB_D_FF_Float_2_9_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder17_Input1_2_0Output, mb_D_FF2_9AugendStage1Output);

    MB_D_FF_Float_2_9_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF2_9AugendStage1Output, mb_D_FF2_9AugendStage2Output);

    Adder_Float_2: entity work.FPAdd_7_24_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF2_9AugendStage2Output, mb_D_FF2_9AddendStage2Output, Adder2_Output_9);

    MB_D_FF_Float_Adder17_Input2_2_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier5_Output_7, mb_D_FFAdder17_Input2_2_0Output);

    MB_D_FF_Float_2_9_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder17_Input2_2_0Output, mb_D_FF2_9AddendStage1Output);

    MB_D_FF_Float_2_9_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF2_9AddendStage1Output, mb_D_FF2_9AddendStage2Output);

    MB_D_FF_Float_Multiplier16_Input1_7_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder2_Output_9, mb_D_FFMultiplier16_Input1_7_0Output);

    MB_D_FF_Float_7_10_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier16_Input1_7_0Output, mb_D_FF7_10MultiplicandStage1Output);

    MB_D_FF_Float_7_10_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF7_10MultiplicandStage1Output, mb_D_FF7_10MultiplicandStage2Output);

    Multiplier_Float_7: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF7_10MultiplicandStage2Output, mb_D_FF7_10MultiplierStage2Output, Multiplier7_Output_10);

    MB_D_FF_Float_Multiplier16_Input2_7_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier4_Output_6, mb_D_FFMultiplier16_Input2_7_0Output);

    MB_D_FF_Float_7_10_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier16_Input2_7_0Output, mb_D_FF7_10MultiplierStage1Output);

    MB_D_FF_Float_7_10_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF7_10MultiplierStage1Output, mb_D_FF7_10MultiplierStage2Output);

    MBRightSHR_Float_8_11: entity work.MBRightSHR(rtl)
    GENERIC MAP (4, NumberOfBits)
    PORT MAP (clk, rst, Multiplier8Weight, mbRightSHR8_11Output);

    MB_D_FF_Float_8_11_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR8_11Output, Multiplier8WeightOutput);

    InputIEEE_Float_8_11: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier8WeightOutput, flopocoMultiplier8WeightOutput);

    MB_D_FF_Float_8_11_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier8WeightOutput, flopocoMultiplier8WeightInput);

    Multiplier_Float_8: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier8WeightInput, mb_D_FF8_11MultiplierStage2Output, Multiplier8_Output_11);

    MB_D_FF_Float_Multiplier20_8_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier20_8_0Input, mb_D_FFMultiplier20_8_0Output);

    MB_D_FF_Float_8_11_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier20_8_0Output, mb_D_FF8_11MultiplierStage1Output);

    MB_D_FF_Float_8_11_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF8_11MultiplierStage1Output, mb_D_FF8_11MultiplierStage2Output);

    MBRightSHR_Float_9_12: entity work.MBRightSHR(rtl)
    GENERIC MAP (4, NumberOfBits)
    PORT MAP (clk, rst, Multiplier9Weight, mbRightSHR9_12Output);

    MB_D_FF_Float_9_12_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR9_12Output, Multiplier9WeightOutput);

    InputIEEE_Float_9_12: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier9WeightOutput, flopocoMultiplier9WeightOutput);

    MB_D_FF_Float_9_12_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier9WeightOutput, flopocoMultiplier9WeightInput);

    Multiplier_Float_9: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier9WeightInput, mb_D_FF9_12MultiplierStage2Output, Multiplier9_Output_12);

    MB_D_FF_Float_Multiplier20_9_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier20_9_0Input, mb_D_FFMultiplier20_9_0Output);

    MB_D_FF_Float_9_12_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier20_9_0Output, mb_D_FF9_12MultiplierStage1Output);

    MB_D_FF_Float_9_12_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF9_12MultiplierStage1Output, mb_D_FF9_12MultiplierStage2Output);

    MB_D_FF_Float_Adder19_Input1_3_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier9_Output_12, mb_D_FFAdder19_Input1_3_0Output);

    MB_D_FF_Float_3_13_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder19_Input1_3_0Output, mb_D_FF3_13AugendStage1Output);

    MB_D_FF_Float_3_13_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF3_13AugendStage1Output, mb_D_FF3_13AugendStage2Output);

    Adder_Float_3: entity work.FPAdd_7_24_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF3_13AugendStage2Output, mb_D_FF3_13AddendStage2Output, Adder3_Output_13);

    MB_D_FF_Float_Adder19_Input2_3_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier8_Output_11, mb_D_FFAdder19_Input2_3_0Output);

    MB_D_FF_Float_3_13_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder19_Input2_3_0Output, mb_D_FF3_13AddendStage1Output);

    MB_D_FF_Float_3_13_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF3_13AddendStage1Output, mb_D_FF3_13AddendStage2Output);

    MB_D_FF_Float_Multiplier18_10_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder3_Output_13, mb_D_FFMultiplier18_10_0Output);

    MB_D_FF_Float_10_14_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier18_10_0Output, mb_D_FF10_14MultiplierStage1Output);

    MB_D_FF_Float_10_14_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF10_14MultiplierStage1Output, mb_D_FF10_14MultiplierStage2Output);

    Multiplier_Float_10: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF10_14MultiplierStage2Output, mb_D_FF10_14MultiplicandStage2Output, Multiplier10_Output_14);

    MBRightSHR_Float_10_14: entity work.MBRightSHR(rtl)
    GENERIC MAP (43, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR10_14Input, mbRightSHR10_14Output);

    MB_D_FF_Float_10_14_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR10_14Output, mb_D_FF10_14MultiplicandStage1Output);

    MB_D_FF_Float_10_14_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF10_14MultiplicandStage1Output, mb_D_FF10_14MultiplicandStage2Output);

    MB_D_FF_Float_Multiplier17_11_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier10_Output_14, mb_D_FFMultiplier17_11_0Output);

    MB_D_FF_Float_11_15_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier17_11_0Output, mb_D_FF11_15MultiplierStage1Output);

    MB_D_FF_Float_11_15_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF11_15MultiplierStage1Output, mb_D_FF11_15MultiplierStage2Output);

    Multiplier_Float_11: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF11_15MultiplierStage2Output, flopocoMultiplier11WeightInput, Multiplier11_Output_15);

    MBRightSHR_Float_11_15: entity work.MBRightSHR(rtl)
    GENERIC MAP (55, NumberOfBits)
    PORT MAP (clk, rst, Multiplier11Weight, mbRightSHR11_15Output);

    MB_D_FF_Float_11_15_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR11_15Output, Multiplier11WeightOutput);

    InputIEEE_Float_11_15: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier11WeightOutput, flopocoMultiplier11WeightOutput);

    MB_D_FF_Float_11_15_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier11WeightOutput, flopocoMultiplier11WeightInput);

    MBRightSHR_Float_12_16: entity work.MBRightSHR(rtl)
    GENERIC MAP (4, NumberOfBits)
    PORT MAP (clk, rst, Multiplier12Weight, mbRightSHR12_16Output);

    MB_D_FF_Float_12_16_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR12_16Output, Multiplier12WeightOutput);

    InputIEEE_Float_12_16: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier12WeightOutput, flopocoMultiplier12WeightOutput);

    MB_D_FF_Float_12_16_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier12WeightOutput, flopocoMultiplier12WeightInput);

    Multiplier_Float_12: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier12WeightInput, mb_D_FF12_16MultiplierStage2Output, Multiplier12_Output_16);

    MB_D_FF_Float_Multiplier20_12_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier20_12_0Input, mb_D_FFMultiplier20_12_0Output);

    MB_D_FF_Float_12_16_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier20_12_0Output, mb_D_FF12_16MultiplierStage1Output);

    MB_D_FF_Float_12_16_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF12_16MultiplierStage1Output, mb_D_FF12_16MultiplierStage2Output);

    MBRightSHR_Float_13_17: entity work.MBRightSHR(rtl)
    GENERIC MAP (4, NumberOfBits)
    PORT MAP (clk, rst, Multiplier13Weight, mbRightSHR13_17Output);

    MB_D_FF_Float_13_17_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR13_17Output, Multiplier13WeightOutput);

    InputIEEE_Float_13_17: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier13WeightOutput, flopocoMultiplier13WeightOutput);

    MB_D_FF_Float_13_17_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier13WeightOutput, flopocoMultiplier13WeightInput);

    Multiplier_Float_13: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier13WeightInput, mb_D_FF13_17MultiplierStage2Output, Multiplier13_Output_17);

    MB_D_FF_Float_Multiplier20_13_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier20_13_0Input, mb_D_FFMultiplier20_13_0Output);

    MB_D_FF_Float_13_17_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier20_13_0Output, mb_D_FF13_17MultiplierStage1Output);

    MB_D_FF_Float_13_17_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF13_17MultiplierStage1Output, mb_D_FF13_17MultiplierStage2Output);

    MB_D_FF_Float_Adder19_Input1_4_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier13_Output_17, mb_D_FFAdder19_Input1_4_0Output);

    MB_D_FF_Float_4_18_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder19_Input1_4_0Output, mb_D_FF4_18AugendStage1Output);

    MB_D_FF_Float_4_18_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF4_18AugendStage1Output, mb_D_FF4_18AugendStage2Output);

    Adder_Float_4: entity work.FPAdd_7_24_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF4_18AugendStage2Output, mb_D_FF4_18AddendStage2Output, Adder4_Output_18);

    MB_D_FF_Float_Adder19_Input2_4_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier12_Output_16, mb_D_FFAdder19_Input2_4_0Output);

    MB_D_FF_Float_4_18_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder19_Input2_4_0Output, mb_D_FF4_18AddendStage1Output);

    MB_D_FF_Float_4_18_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF4_18AddendStage1Output, mb_D_FF4_18AddendStage2Output);

    MB_D_FF_Float_Multiplier18_14_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder4_Output_18, mb_D_FFMultiplier18_14_0Output);

    MB_D_FF_Float_14_19_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier18_14_0Output, mb_D_FF14_19MultiplierStage1Output);

    MB_D_FF_Float_14_19_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF14_19MultiplierStage1Output, mb_D_FF14_19MultiplierStage2Output);

    Multiplier_Float_14: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF14_19MultiplierStage2Output, mb_D_FF14_19MultiplicandStage2Output, Multiplier14_Output_19);

    MBRightSHR_Float_14_19: entity work.MBRightSHR(rtl)
    GENERIC MAP (43, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR14_19Input, mbRightSHR14_19Output);

    MB_D_FF_Float_14_19_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR14_19Output, mb_D_FF14_19MultiplicandStage1Output);

    MB_D_FF_Float_14_19_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF14_19MultiplicandStage1Output, mb_D_FF14_19MultiplicandStage2Output);

    MB_D_FF_Float_Multiplier17_15_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier14_Output_19, mb_D_FFMultiplier17_15_0Output);

    MB_D_FF_Float_15_20_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier17_15_0Output, mb_D_FF15_20MultiplierStage1Output);

    MB_D_FF_Float_15_20_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF15_20MultiplierStage1Output, mb_D_FF15_20MultiplierStage2Output);

    Multiplier_Float_15: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF15_20MultiplierStage2Output, flopocoMultiplier15WeightInput, Multiplier15_Output_20);

    MBRightSHR_Float_15_20: entity work.MBRightSHR(rtl)
    GENERIC MAP (55, NumberOfBits)
    PORT MAP (clk, rst, Multiplier15Weight, mbRightSHR15_20Output);

    MB_D_FF_Float_15_20_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR15_20Output, Multiplier15WeightOutput);

    InputIEEE_Float_15_20: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier15WeightOutput, flopocoMultiplier15WeightOutput);

    MB_D_FF_Float_15_20_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier15WeightOutput, flopocoMultiplier15WeightInput);

    MB_D_FF_Float_Adder16_Input1_5_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier15_Output_20, mb_D_FFAdder16_Input1_5_0Output);

    MB_D_FF_Float_5_21_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder16_Input1_5_0Output, mb_D_FF5_21AugendStage1Output);

    MB_D_FF_Float_5_21_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF5_21AugendStage1Output, mb_D_FF5_21AugendStage2Output);

    Adder_Float_5: entity work.FPAdd_7_24_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF5_21AugendStage2Output, mb_D_FF5_21AddendStage2Output, Adder5_Output_21);

    MB_D_FF_Float_Adder16_Input2_5_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier11_Output_15, mb_D_FFAdder16_Input2_5_0Output);

    MB_D_FF_Float_5_21_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder16_Input2_5_0Output, mb_D_FF5_21AddendStage1Output);

    MB_D_FF_Float_5_21_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF5_21AddendStage1Output, mb_D_FF5_21AddendStage2Output);

    MB_D_FF_Float_Multiplier15_Input1_16_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder5_Output_21, mb_D_FFMultiplier15_Input1_16_0Output);

    MB_D_FF_Float_16_22_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier15_Input1_16_0Output, mb_D_FF16_22MultiplicandStage1Output);

    MB_D_FF_Float_16_22_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF16_22MultiplicandStage1Output, mb_D_FF16_22MultiplicandStage2Output);

    Multiplier_Float_16: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF16_22MultiplicandStage2Output, mb_D_FF16_22MultiplierStage2Output, Multiplier16_Output_22);

    MB_D_FF_Float_Multiplier15_Input2_16_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier7_Output_10, mb_D_FFMultiplier15_Input2_16_0Output);

    MB_D_FF_Float_16_22_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier15_Input2_16_0Output, mb_D_FF16_22MultiplierStage1Output);

    MB_D_FF_Float_16_22_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF16_22MultiplierStage1Output, mb_D_FF16_22MultiplierStage2Output);

    MBRightSHR_Float_17_Input123: entity work.MBRightSHR(rtl)
    GENERIC MAP (67, NumberOfBits)
    PORT MAP (clk, rst, Multiplier17Weight, mbRightSHR17_Input1_23Output);

    MB_D_FF_Float_17_23_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR17_Input1_23Output, Multiplier17WeightOutput);

    InputIEEE_Float_17_23: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier17WeightOutput, flopocoMultiplier17WeightOutput);

    MB_D_FF_Float_17_23_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier17WeightOutput, flopocoMultiplier17WeightInput);

    Multiplier_Float_17: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier17WeightInput, mb_D_FF17_23MultiplierStage2Output, Multiplier17_Output_23);

    MBRightSHR_Float_17_Input2_23: entity work.MBRightSHR(rtl)
    GENERIC MAP (67, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR17_Input2_23Input, mbRightSHR17_Input2_23Output);

    MB_D_FF_Float_17_23_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR17_Input2_23Output, mb_D_FF17_23MultiplierStage1Output);

    MB_D_FF_Float_17_23_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF17_23MultiplierStage1Output, mb_D_FF17_23MultiplierStage2Output);

    MBRightSHR_Float_18_Input124: entity work.MBRightSHR(rtl)
    GENERIC MAP (67, NumberOfBits)
    PORT MAP (clk, rst, Multiplier18Weight, mbRightSHR18_Input1_24Output);

    MB_D_FF_Float_18_24_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR18_Input1_24Output, Multiplier18WeightOutput);

    InputIEEE_Float_18_24: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier18WeightOutput, flopocoMultiplier18WeightOutput);

    MB_D_FF_Float_18_24_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier18WeightOutput, flopocoMultiplier18WeightInput);

    Multiplier_Float_18: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier18WeightInput, mb_D_FF18_24MultiplierStage2Output, Multiplier18_Output_24);

    MBRightSHR_Float_18_Input2_24: entity work.MBRightSHR(rtl)
    GENERIC MAP (67, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR18_Input2_24Input, mbRightSHR18_Input2_24Output);

    MB_D_FF_Float_18_24_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR18_Input2_24Output, mb_D_FF18_24MultiplierStage1Output);

    MB_D_FF_Float_18_24_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF18_24MultiplierStage1Output, mb_D_FF18_24MultiplierStage2Output);

    MB_D_FF_Float_Adder15_Input1_6_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier18_Output_24, mb_D_FFAdder15_Input1_6_0Output);

    MB_D_FF_Float_6_25_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder15_Input1_6_0Output, mb_D_FF6_25AugendStage1Output);

    MB_D_FF_Float_6_25_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF6_25AugendStage1Output, mb_D_FF6_25AugendStage2Output);

    Adder_Float_6: entity work.FPAdd_7_24_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF6_25AugendStage2Output, mb_D_FF6_25AddendStage2Output, Adder6_Output_25);

    MB_D_FF_Float_Adder15_Input2_6_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier17_Output_23, mb_D_FFAdder15_Input2_6_0Output);

    MB_D_FF_Float_6_25_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder15_Input2_6_0Output, mb_D_FF6_25AddendStage1Output);

    MB_D_FF_Float_6_25_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF6_25AddendStage1Output, mb_D_FF6_25AddendStage2Output);

    MB_D_FF_Float_Multiplier14_Input1_19_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder6_Output_25, mb_D_FFMultiplier14_Input1_19_0Output);

    MB_D_FF_Float_19_26_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier14_Input1_19_0Output, mb_D_FF19_26MultiplicandStage1Output);

    MB_D_FF_Float_19_26_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF19_26MultiplicandStage1Output, mb_D_FF19_26MultiplicandStage2Output);

    Multiplier_Float_19: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF19_26MultiplicandStage2Output, mb_D_FF19_26MultiplierStage2Output, Multiplier19_Output_26);

    MB_D_FF_Float_Multiplier14_Input2_19_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier16_Output_22, mb_D_FFMultiplier14_Input2_19_0Output);

    MB_D_FF_Float_19_26_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier14_Input2_19_0Output, mb_D_FF19_26MultiplierStage1Output);

    MB_D_FF_Float_19_26_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF19_26MultiplierStage1Output, mb_D_FF19_26MultiplierStage2Output);

    MBRightSHR_Float_20_Input127: entity work.MBRightSHR(rtl)
    GENERIC MAP (94, NumberOfBits)
    PORT MAP (clk, rst, Multiplier20Weight, mbRightSHR20_Input1_27Output);

    MB_D_FF_Float_20_27_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR20_Input1_27Output, Multiplier20WeightOutput);

    InputIEEE_Float_20_27: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier20WeightOutput, flopocoMultiplier20WeightOutput);

    MB_D_FF_Float_20_27_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier20WeightOutput, flopocoMultiplier20WeightInput);

    Multiplier_Float_20: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier20WeightInput, mb_D_FF20_27MultiplierStage2Output, Multiplier20_Output_27);

    MBRightSHR_Float_20_Input2_27: entity work.MBRightSHR(rtl)
    GENERIC MAP (94, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR20_Input2_27Input, mbRightSHR20_Input2_27Output);

    MB_D_FF_Float_20_27_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR20_Input2_27Output, mb_D_FF20_27MultiplierStage1Output);

    MB_D_FF_Float_20_27_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF20_27MultiplierStage1Output, mb_D_FF20_27MultiplierStage2Output);

    MBRightSHR_Float_21_Input128: entity work.MBRightSHR(rtl)
    GENERIC MAP (94, NumberOfBits)
    PORT MAP (clk, rst, Multiplier21Weight, mbRightSHR21_Input1_28Output);

    MB_D_FF_Float_21_28_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR21_Input1_28Output, Multiplier21WeightOutput);

    InputIEEE_Float_21_28: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier21WeightOutput, flopocoMultiplier21WeightOutput);

    MB_D_FF_Float_21_28_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier21WeightOutput, flopocoMultiplier21WeightInput);

    Multiplier_Float_21: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier21WeightInput, mb_D_FF21_28MultiplierStage2Output, Multiplier21_Output_28);

    MBRightSHR_Float_21_Input2_28: entity work.MBRightSHR(rtl)
    GENERIC MAP (94, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR21_Input2_28Input, mbRightSHR21_Input2_28Output);

    MB_D_FF_Float_21_28_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR21_Input2_28Output, mb_D_FF21_28MultiplierStage1Output);

    MB_D_FF_Float_21_28_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF21_28MultiplierStage1Output, mb_D_FF21_28MultiplierStage2Output);

    MB_D_FF_Float_Adder14_Input1_7_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier21_Output_28, mb_D_FFAdder14_Input1_7_0Output);

    MB_D_FF_Float_7_29_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder14_Input1_7_0Output, mb_D_FF7_29AugendStage1Output);

    MB_D_FF_Float_7_29_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF7_29AugendStage1Output, mb_D_FF7_29AugendStage2Output);

    Adder_Float_7: entity work.FPAdd_7_24_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF7_29AugendStage2Output, mb_D_FF7_29AddendStage2Output, Adder7_Output_29);

    MB_D_FF_Float_Adder14_Input2_7_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier20_Output_27, mb_D_FFAdder14_Input2_7_0Output);

    MB_D_FF_Float_7_29_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder14_Input2_7_0Output, mb_D_FF7_29AddendStage1Output);

    MB_D_FF_Float_7_29_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF7_29AddendStage1Output, mb_D_FF7_29AddendStage2Output);

    MB_D_FF_Float_Multiplier13_Input1_22_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder7_Output_29, mb_D_FFMultiplier13_Input1_22_0Output);

    MB_D_FF_Float_22_30_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier13_Input1_22_0Output, mb_D_FF22_30MultiplicandStage1Output);

    MB_D_FF_Float_22_30_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF22_30MultiplicandStage1Output, mb_D_FF22_30MultiplicandStage2Output);

    Multiplier_Float_22: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF22_30MultiplicandStage2Output, mb_D_FF22_30MultiplierStage2Output, Multiplier22_Output_30);

    MB_D_FF_Float_Multiplier13_Input2_22_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier19_Output_26, mb_D_FFMultiplier13_Input2_22_0Output);

    MB_D_FF_Float_22_30_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier13_Input2_22_0Output, mb_D_FF22_30MultiplierStage1Output);

    MB_D_FF_Float_22_30_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF22_30MultiplierStage1Output, mb_D_FF22_30MultiplierStage2Output);

    MBRightSHR_Float_23_Input131: entity work.MBRightSHR(rtl)
    GENERIC MAP (106, NumberOfBits)
    PORT MAP (clk, rst, Multiplier23Weight, mbRightSHR23_Input1_31Output);

    MB_D_FF_Float_23_31_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR23_Input1_31Output, Multiplier23WeightOutput);

    InputIEEE_Float_23_31: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier23WeightOutput, flopocoMultiplier23WeightOutput);

    MB_D_FF_Float_23_31_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier23WeightOutput, flopocoMultiplier23WeightInput);

    Multiplier_Float_23: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier23WeightInput, mb_D_FF23_31MultiplierStage2Output, Multiplier23_Output_31);

    MBRightSHR_Float_23_Input2_31: entity work.MBRightSHR(rtl)
    GENERIC MAP (106, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR23_Input2_31Input, mbRightSHR23_Input2_31Output);

    MB_D_FF_Float_23_31_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR23_Input2_31Output, mb_D_FF23_31MultiplierStage1Output);

    MB_D_FF_Float_23_31_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF23_31MultiplierStage1Output, mb_D_FF23_31MultiplierStage2Output);

    MBRightSHR_Float_24_Input132: entity work.MBRightSHR(rtl)
    GENERIC MAP (106, NumberOfBits)
    PORT MAP (clk, rst, Multiplier24Weight, mbRightSHR24_Input1_32Output);

    MB_D_FF_Float_24_32_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR24_Input1_32Output, Multiplier24WeightOutput);

    InputIEEE_Float_24_32: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier24WeightOutput, flopocoMultiplier24WeightOutput);

    MB_D_FF_Float_24_32_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier24WeightOutput, flopocoMultiplier24WeightInput);

    Multiplier_Float_24: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier24WeightInput, mb_D_FF24_32MultiplierStage2Output, Multiplier24_Output_32);

    MBRightSHR_Float_24_Input2_32: entity work.MBRightSHR(rtl)
    GENERIC MAP (106, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR24_Input2_32Input, mbRightSHR24_Input2_32Output);

    MB_D_FF_Float_24_32_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR24_Input2_32Output, mb_D_FF24_32MultiplierStage1Output);

    MB_D_FF_Float_24_32_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF24_32MultiplierStage1Output, mb_D_FF24_32MultiplierStage2Output);

    MB_D_FF_Float_Adder13_Input1_8_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier24_Output_32, mb_D_FFAdder13_Input1_8_0Output);

    MB_D_FF_Float_8_33_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder13_Input1_8_0Output, mb_D_FF8_33AugendStage1Output);

    MB_D_FF_Float_8_33_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF8_33AugendStage1Output, mb_D_FF8_33AugendStage2Output);

    Adder_Float_8: entity work.FPAdd_7_24_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF8_33AugendStage2Output, mb_D_FF8_33AddendStage2Output, Adder8_Output_33);

    MB_D_FF_Float_Adder13_Input2_8_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier23_Output_31, mb_D_FFAdder13_Input2_8_0Output);

    MB_D_FF_Float_8_33_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder13_Input2_8_0Output, mb_D_FF8_33AddendStage1Output);

    MB_D_FF_Float_8_33_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF8_33AddendStage1Output, mb_D_FF8_33AddendStage2Output);

    MB_D_FF_Float_Multiplier12_Input1_25_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder8_Output_33, mb_D_FFMultiplier12_Input1_25_0Output);

    MB_D_FF_Float_25_34_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier12_Input1_25_0Output, mb_D_FF25_34MultiplicandStage1Output);

    MB_D_FF_Float_25_34_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF25_34MultiplicandStage1Output, mb_D_FF25_34MultiplicandStage2Output);

    Multiplier_Float_25: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF25_34MultiplicandStage2Output, mb_D_FF25_34MultiplierStage2Output, Multiplier25_Output_34);

    MB_D_FF_Float_Multiplier12_Input2_25_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier22_Output_30, mb_D_FFMultiplier12_Input2_25_0Output);

    MB_D_FF_Float_25_34_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier12_Input2_25_0Output, mb_D_FF25_34MultiplierStage1Output);

    MB_D_FF_Float_25_34_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF25_34MultiplierStage1Output, mb_D_FF25_34MultiplierStage2Output);

    MBRightSHR_Float_26_Input135: entity work.MBRightSHR(rtl)
    GENERIC MAP (118, NumberOfBits)
    PORT MAP (clk, rst, Multiplier26Weight, mbRightSHR26_Input1_35Output);

    MB_D_FF_Float_26_35_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR26_Input1_35Output, Multiplier26WeightOutput);

    InputIEEE_Float_26_35: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier26WeightOutput, flopocoMultiplier26WeightOutput);

    MB_D_FF_Float_26_35_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier26WeightOutput, flopocoMultiplier26WeightInput);

    Multiplier_Float_26: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier26WeightInput, mb_D_FF26_35MultiplierStage2Output, Multiplier26_Output_35);

    MBRightSHR_Float_26_Input2_35: entity work.MBRightSHR(rtl)
    GENERIC MAP (118, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR26_Input2_35Input, mbRightSHR26_Input2_35Output);

    MB_D_FF_Float_26_35_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR26_Input2_35Output, mb_D_FF26_35MultiplierStage1Output);

    MB_D_FF_Float_26_35_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF26_35MultiplierStage1Output, mb_D_FF26_35MultiplierStage2Output);

    MBRightSHR_Float_27_Input136: entity work.MBRightSHR(rtl)
    GENERIC MAP (118, NumberOfBits)
    PORT MAP (clk, rst, Multiplier27Weight, mbRightSHR27_Input1_36Output);

    MB_D_FF_Float_27_36_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR27_Input1_36Output, Multiplier27WeightOutput);

    InputIEEE_Float_27_36: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier27WeightOutput, flopocoMultiplier27WeightOutput);

    MB_D_FF_Float_27_36_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier27WeightOutput, flopocoMultiplier27WeightInput);

    Multiplier_Float_27: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier27WeightInput, mb_D_FF27_36MultiplierStage2Output, Multiplier27_Output_36);

    MBRightSHR_Float_27_Input2_36: entity work.MBRightSHR(rtl)
    GENERIC MAP (118, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR27_Input2_36Input, mbRightSHR27_Input2_36Output);

    MB_D_FF_Float_27_36_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR27_Input2_36Output, mb_D_FF27_36MultiplierStage1Output);

    MB_D_FF_Float_27_36_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF27_36MultiplierStage1Output, mb_D_FF27_36MultiplierStage2Output);

    MB_D_FF_Float_Adder12_Input1_9_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier27_Output_36, mb_D_FFAdder12_Input1_9_0Output);

    MB_D_FF_Float_9_37_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder12_Input1_9_0Output, mb_D_FF9_37AugendStage1Output);

    MB_D_FF_Float_9_37_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF9_37AugendStage1Output, mb_D_FF9_37AugendStage2Output);

    Adder_Float_9: entity work.FPAdd_7_24_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF9_37AugendStage2Output, mb_D_FF9_37AddendStage2Output, Adder9_Output_37);

    MB_D_FF_Float_Adder12_Input2_9_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier26_Output_35, mb_D_FFAdder12_Input2_9_0Output);

    MB_D_FF_Float_9_37_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder12_Input2_9_0Output, mb_D_FF9_37AddendStage1Output);

    MB_D_FF_Float_9_37_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF9_37AddendStage1Output, mb_D_FF9_37AddendStage2Output);

    MB_D_FF_Float_Multiplier11_Input1_28_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder9_Output_37, mb_D_FFMultiplier11_Input1_28_0Output);

    MB_D_FF_Float_28_38_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier11_Input1_28_0Output, mb_D_FF28_38MultiplicandStage1Output);

    MB_D_FF_Float_28_38_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF28_38MultiplicandStage1Output, mb_D_FF28_38MultiplicandStage2Output);

    Multiplier_Float_28: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF28_38MultiplicandStage2Output, mb_D_FF28_38MultiplierStage2Output, Multiplier28_Output_38);

    MB_D_FF_Float_Multiplier11_Input2_28_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier25_Output_34, mb_D_FFMultiplier11_Input2_28_0Output);

    MB_D_FF_Float_28_38_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier11_Input2_28_0Output, mb_D_FF28_38MultiplierStage1Output);

    MB_D_FF_Float_28_38_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF28_38MultiplierStage1Output, mb_D_FF28_38MultiplierStage2Output);

    MBRightSHR_Float_29_Input139: entity work.MBRightSHR(rtl)
    GENERIC MAP (130, NumberOfBits)
    PORT MAP (clk, rst, Multiplier29Weight, mbRightSHR29_Input1_39Output);

    MB_D_FF_Float_29_39_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR29_Input1_39Output, Multiplier29WeightOutput);

    InputIEEE_Float_29_39: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier29WeightOutput, flopocoMultiplier29WeightOutput);

    MB_D_FF_Float_29_39_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier29WeightOutput, flopocoMultiplier29WeightInput);

    Multiplier_Float_29: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier29WeightInput, mb_D_FF29_39MultiplierStage2Output, Multiplier29_Output_39);

    MBRightSHR_Float_29_Input2_39: entity work.MBRightSHR(rtl)
    GENERIC MAP (130, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR29_Input2_39Input, mbRightSHR29_Input2_39Output);

    MB_D_FF_Float_29_39_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR29_Input2_39Output, mb_D_FF29_39MultiplierStage1Output);

    MB_D_FF_Float_29_39_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF29_39MultiplierStage1Output, mb_D_FF29_39MultiplierStage2Output);

    MBRightSHR_Float_30_Input140: entity work.MBRightSHR(rtl)
    GENERIC MAP (130, NumberOfBits)
    PORT MAP (clk, rst, Multiplier30Weight, mbRightSHR30_Input1_40Output);

    MB_D_FF_Float_30_40_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR30_Input1_40Output, Multiplier30WeightOutput);

    InputIEEE_Float_30_40: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier30WeightOutput, flopocoMultiplier30WeightOutput);

    MB_D_FF_Float_30_40_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier30WeightOutput, flopocoMultiplier30WeightInput);

    Multiplier_Float_30: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier30WeightInput, mb_D_FF30_40MultiplierStage2Output, Multiplier30_Output_40);

    MBRightSHR_Float_30_Input2_40: entity work.MBRightSHR(rtl)
    GENERIC MAP (130, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR30_Input2_40Input, mbRightSHR30_Input2_40Output);

    MB_D_FF_Float_30_40_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR30_Input2_40Output, mb_D_FF30_40MultiplierStage1Output);

    MB_D_FF_Float_30_40_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF30_40MultiplierStage1Output, mb_D_FF30_40MultiplierStage2Output);

    MB_D_FF_Float_Adder11_Input1_10_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier30_Output_40, mb_D_FFAdder11_Input1_10_0Output);

    MB_D_FF_Float_10_41_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder11_Input1_10_0Output, mb_D_FF10_41AugendStage1Output);

    MB_D_FF_Float_10_41_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF10_41AugendStage1Output, mb_D_FF10_41AugendStage2Output);

    Adder_Float_10: entity work.FPAdd_7_24_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF10_41AugendStage2Output, mb_D_FF10_41AddendStage2Output, Adder10_Output_41);

    MB_D_FF_Float_Adder11_Input2_10_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier29_Output_39, mb_D_FFAdder11_Input2_10_0Output);

    MB_D_FF_Float_10_41_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder11_Input2_10_0Output, mb_D_FF10_41AddendStage1Output);

    MB_D_FF_Float_10_41_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF10_41AddendStage1Output, mb_D_FF10_41AddendStage2Output);

    MB_D_FF_Float_Multiplier10_Input1_31_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder10_Output_41, mb_D_FFMultiplier10_Input1_31_0Output);

    MB_D_FF_Float_31_42_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier10_Input1_31_0Output, mb_D_FF31_42MultiplicandStage1Output);

    MB_D_FF_Float_31_42_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF31_42MultiplicandStage1Output, mb_D_FF31_42MultiplicandStage2Output);

    Multiplier_Float_31: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF31_42MultiplicandStage2Output, mb_D_FF31_42MultiplierStage2Output, Multiplier31_Output_42);

    MB_D_FF_Float_Multiplier10_Input2_31_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier28_Output_38, mb_D_FFMultiplier10_Input2_31_0Output);

    MB_D_FF_Float_31_42_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier10_Input2_31_0Output, mb_D_FF31_42MultiplierStage1Output);

    MB_D_FF_Float_31_42_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF31_42MultiplierStage1Output, mb_D_FF31_42MultiplierStage2Output);

    MBRightSHR_Float_32_Input143: entity work.MBRightSHR(rtl)
    GENERIC MAP (142, NumberOfBits)
    PORT MAP (clk, rst, Multiplier32Weight, mbRightSHR32_Input1_43Output);

    MB_D_FF_Float_32_43_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR32_Input1_43Output, Multiplier32WeightOutput);

    InputIEEE_Float_32_43: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier32WeightOutput, flopocoMultiplier32WeightOutput);

    MB_D_FF_Float_32_43_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier32WeightOutput, flopocoMultiplier32WeightInput);

    Multiplier_Float_32: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier32WeightInput, mb_D_FF32_43MultiplierStage2Output, Multiplier32_Output_43);

    MBRightSHR_Float_32_Input2_43: entity work.MBRightSHR(rtl)
    GENERIC MAP (142, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR32_Input2_43Input, mbRightSHR32_Input2_43Output);

    MB_D_FF_Float_32_43_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR32_Input2_43Output, mb_D_FF32_43MultiplierStage1Output);

    MB_D_FF_Float_32_43_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF32_43MultiplierStage1Output, mb_D_FF32_43MultiplierStage2Output);

    MBRightSHR_Float_33_Input144: entity work.MBRightSHR(rtl)
    GENERIC MAP (142, NumberOfBits)
    PORT MAP (clk, rst, Multiplier33Weight, mbRightSHR33_Input1_44Output);

    MB_D_FF_Float_33_44_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR33_Input1_44Output, Multiplier33WeightOutput);

    InputIEEE_Float_33_44: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier33WeightOutput, flopocoMultiplier33WeightOutput);

    MB_D_FF_Float_33_44_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier33WeightOutput, flopocoMultiplier33WeightInput);

    Multiplier_Float_33: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier33WeightInput, mb_D_FF33_44MultiplierStage2Output, Multiplier33_Output_44);

    MBRightSHR_Float_33_Input2_44: entity work.MBRightSHR(rtl)
    GENERIC MAP (142, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR33_Input2_44Input, mbRightSHR33_Input2_44Output);

    MB_D_FF_Float_33_44_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR33_Input2_44Output, mb_D_FF33_44MultiplierStage1Output);

    MB_D_FF_Float_33_44_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF33_44MultiplierStage1Output, mb_D_FF33_44MultiplierStage2Output);

    MB_D_FF_Float_Adder10_Input1_11_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier33_Output_44, mb_D_FFAdder10_Input1_11_0Output);

    MB_D_FF_Float_11_45_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder10_Input1_11_0Output, mb_D_FF11_45AugendStage1Output);

    MB_D_FF_Float_11_45_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF11_45AugendStage1Output, mb_D_FF11_45AugendStage2Output);

    Adder_Float_11: entity work.FPAdd_7_24_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF11_45AugendStage2Output, mb_D_FF11_45AddendStage2Output, Adder11_Output_45);

    MB_D_FF_Float_Adder10_Input2_11_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier32_Output_43, mb_D_FFAdder10_Input2_11_0Output);

    MB_D_FF_Float_11_45_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder10_Input2_11_0Output, mb_D_FF11_45AddendStage1Output);

    MB_D_FF_Float_11_45_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF11_45AddendStage1Output, mb_D_FF11_45AddendStage2Output);

    MB_D_FF_Float_Multiplier9_Input1_34_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder11_Output_45, mb_D_FFMultiplier9_Input1_34_0Output);

    MB_D_FF_Float_34_46_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier9_Input1_34_0Output, mb_D_FF34_46MultiplicandStage1Output);

    MB_D_FF_Float_34_46_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF34_46MultiplicandStage1Output, mb_D_FF34_46MultiplicandStage2Output);

    Multiplier_Float_34: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF34_46MultiplicandStage2Output, mb_D_FF34_46MultiplierStage2Output, Multiplier34_Output_46);

    MB_D_FF_Float_Multiplier9_Input2_34_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier31_Output_42, mb_D_FFMultiplier9_Input2_34_0Output);

    MB_D_FF_Float_34_46_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier9_Input2_34_0Output, mb_D_FF34_46MultiplierStage1Output);

    MB_D_FF_Float_34_46_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF34_46MultiplierStage1Output, mb_D_FF34_46MultiplierStage2Output);

    MBRightSHR_Float_35_Input147: entity work.MBRightSHR(rtl)
    GENERIC MAP (154, NumberOfBits)
    PORT MAP (clk, rst, Multiplier35Weight, mbRightSHR35_Input1_47Output);

    MB_D_FF_Float_35_47_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR35_Input1_47Output, Multiplier35WeightOutput);

    InputIEEE_Float_35_47: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier35WeightOutput, flopocoMultiplier35WeightOutput);

    MB_D_FF_Float_35_47_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier35WeightOutput, flopocoMultiplier35WeightInput);

    Multiplier_Float_35: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier35WeightInput, mb_D_FF35_47MultiplierStage2Output, Multiplier35_Output_47);

    MBRightSHR_Float_35_Input2_47: entity work.MBRightSHR(rtl)
    GENERIC MAP (154, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR35_Input2_47Input, mbRightSHR35_Input2_47Output);

    MB_D_FF_Float_35_47_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR35_Input2_47Output, mb_D_FF35_47MultiplierStage1Output);

    MB_D_FF_Float_35_47_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF35_47MultiplierStage1Output, mb_D_FF35_47MultiplierStage2Output);

    MBRightSHR_Float_36_Input148: entity work.MBRightSHR(rtl)
    GENERIC MAP (154, NumberOfBits)
    PORT MAP (clk, rst, Multiplier36Weight, mbRightSHR36_Input1_48Output);

    MB_D_FF_Float_36_48_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR36_Input1_48Output, Multiplier36WeightOutput);

    InputIEEE_Float_36_48: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier36WeightOutput, flopocoMultiplier36WeightOutput);

    MB_D_FF_Float_36_48_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier36WeightOutput, flopocoMultiplier36WeightInput);

    Multiplier_Float_36: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier36WeightInput, mb_D_FF36_48MultiplierStage2Output, Multiplier36_Output_48);

    MBRightSHR_Float_36_Input2_48: entity work.MBRightSHR(rtl)
    GENERIC MAP (154, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR36_Input2_48Input, mbRightSHR36_Input2_48Output);

    MB_D_FF_Float_36_48_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR36_Input2_48Output, mb_D_FF36_48MultiplierStage1Output);

    MB_D_FF_Float_36_48_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF36_48MultiplierStage1Output, mb_D_FF36_48MultiplierStage2Output);

    MB_D_FF_Float_Adder9_Input1_12_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier36_Output_48, mb_D_FFAdder9_Input1_12_0Output);

    MB_D_FF_Float_12_49_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder9_Input1_12_0Output, mb_D_FF12_49AugendStage1Output);

    MB_D_FF_Float_12_49_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF12_49AugendStage1Output, mb_D_FF12_49AugendStage2Output);

    Adder_Float_12: entity work.FPAdd_7_24_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF12_49AugendStage2Output, mb_D_FF12_49AddendStage2Output, Adder12_Output_49);

    MB_D_FF_Float_Adder9_Input2_12_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier35_Output_47, mb_D_FFAdder9_Input2_12_0Output);

    MB_D_FF_Float_12_49_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder9_Input2_12_0Output, mb_D_FF12_49AddendStage1Output);

    MB_D_FF_Float_12_49_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF12_49AddendStage1Output, mb_D_FF12_49AddendStage2Output);

    MB_D_FF_Float_Multiplier8_Input1_37_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder12_Output_49, mb_D_FFMultiplier8_Input1_37_0Output);

    MB_D_FF_Float_37_50_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier8_Input1_37_0Output, mb_D_FF37_50MultiplicandStage1Output);

    MB_D_FF_Float_37_50_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF37_50MultiplicandStage1Output, mb_D_FF37_50MultiplicandStage2Output);

    Multiplier_Float_37: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF37_50MultiplicandStage2Output, mb_D_FF37_50MultiplierStage2Output, Multiplier37_Output_50);

    MB_D_FF_Float_Multiplier8_Input2_37_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier34_Output_46, mb_D_FFMultiplier8_Input2_37_0Output);

    MB_D_FF_Float_37_50_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier8_Input2_37_0Output, mb_D_FF37_50MultiplierStage1Output);

    MB_D_FF_Float_37_50_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF37_50MultiplierStage1Output, mb_D_FF37_50MultiplierStage2Output);

    MBRightSHR_Float_38_Input151: entity work.MBRightSHR(rtl)
    GENERIC MAP (166, NumberOfBits)
    PORT MAP (clk, rst, Multiplier38Weight, mbRightSHR38_Input1_51Output);

    MB_D_FF_Float_38_51_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR38_Input1_51Output, Multiplier38WeightOutput);

    InputIEEE_Float_38_51: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier38WeightOutput, flopocoMultiplier38WeightOutput);

    MB_D_FF_Float_38_51_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier38WeightOutput, flopocoMultiplier38WeightInput);

    Multiplier_Float_38: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier38WeightInput, mb_D_FF38_51MultiplierStage2Output, Multiplier38_Output_51);

    MBRightSHR_Float_38_Input2_51: entity work.MBRightSHR(rtl)
    GENERIC MAP (166, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR38_Input2_51Input, mbRightSHR38_Input2_51Output);

    MB_D_FF_Float_38_51_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR38_Input2_51Output, mb_D_FF38_51MultiplierStage1Output);

    MB_D_FF_Float_38_51_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF38_51MultiplierStage1Output, mb_D_FF38_51MultiplierStage2Output);

    MBRightSHR_Float_39_Input152: entity work.MBRightSHR(rtl)
    GENERIC MAP (166, NumberOfBits)
    PORT MAP (clk, rst, Multiplier39Weight, mbRightSHR39_Input1_52Output);

    MB_D_FF_Float_39_52_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR39_Input1_52Output, Multiplier39WeightOutput);

    InputIEEE_Float_39_52: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier39WeightOutput, flopocoMultiplier39WeightOutput);

    MB_D_FF_Float_39_52_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier39WeightOutput, flopocoMultiplier39WeightInput);

    Multiplier_Float_39: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier39WeightInput, mb_D_FF39_52MultiplierStage2Output, Multiplier39_Output_52);

    MBRightSHR_Float_39_Input2_52: entity work.MBRightSHR(rtl)
    GENERIC MAP (166, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR39_Input2_52Input, mbRightSHR39_Input2_52Output);

    MB_D_FF_Float_39_52_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR39_Input2_52Output, mb_D_FF39_52MultiplierStage1Output);

    MB_D_FF_Float_39_52_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF39_52MultiplierStage1Output, mb_D_FF39_52MultiplierStage2Output);

    MB_D_FF_Float_Adder8_Input1_13_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier39_Output_52, mb_D_FFAdder8_Input1_13_0Output);

    MB_D_FF_Float_13_53_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder8_Input1_13_0Output, mb_D_FF13_53AugendStage1Output);

    MB_D_FF_Float_13_53_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF13_53AugendStage1Output, mb_D_FF13_53AugendStage2Output);

    Adder_Float_13: entity work.FPAdd_7_24_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF13_53AugendStage2Output, mb_D_FF13_53AddendStage2Output, Adder13_Output_53);

    MB_D_FF_Float_Adder8_Input2_13_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier38_Output_51, mb_D_FFAdder8_Input2_13_0Output);

    MB_D_FF_Float_13_53_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder8_Input2_13_0Output, mb_D_FF13_53AddendStage1Output);

    MB_D_FF_Float_13_53_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF13_53AddendStage1Output, mb_D_FF13_53AddendStage2Output);

    MB_D_FF_Float_Multiplier7_Input1_40_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder13_Output_53, mb_D_FFMultiplier7_Input1_40_0Output);

    MB_D_FF_Float_40_54_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier7_Input1_40_0Output, mb_D_FF40_54MultiplicandStage1Output);

    MB_D_FF_Float_40_54_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF40_54MultiplicandStage1Output, mb_D_FF40_54MultiplicandStage2Output);

    Multiplier_Float_40: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF40_54MultiplicandStage2Output, mb_D_FF40_54MultiplierStage2Output, Multiplier40_Output_54);

    MB_D_FF_Float_Multiplier7_Input2_40_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier37_Output_50, mb_D_FFMultiplier7_Input2_40_0Output);

    MB_D_FF_Float_40_54_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier7_Input2_40_0Output, mb_D_FF40_54MultiplierStage1Output);

    MB_D_FF_Float_40_54_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF40_54MultiplierStage1Output, mb_D_FF40_54MultiplierStage2Output);

    MBRightSHR_Float_41_Input155: entity work.MBRightSHR(rtl)
    GENERIC MAP (178, NumberOfBits)
    PORT MAP (clk, rst, Multiplier41Weight, mbRightSHR41_Input1_55Output);

    MB_D_FF_Float_41_55_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR41_Input1_55Output, Multiplier41WeightOutput);

    InputIEEE_Float_41_55: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier41WeightOutput, flopocoMultiplier41WeightOutput);

    MB_D_FF_Float_41_55_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier41WeightOutput, flopocoMultiplier41WeightInput);

    Multiplier_Float_41: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier41WeightInput, mb_D_FF41_55MultiplierStage2Output, Multiplier41_Output_55);

    MBRightSHR_Float_41_Input2_55: entity work.MBRightSHR(rtl)
    GENERIC MAP (178, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR41_Input2_55Input, mbRightSHR41_Input2_55Output);

    MB_D_FF_Float_41_55_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR41_Input2_55Output, mb_D_FF41_55MultiplierStage1Output);

    MB_D_FF_Float_41_55_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF41_55MultiplierStage1Output, mb_D_FF41_55MultiplierStage2Output);

    MBRightSHR_Float_42_Input156: entity work.MBRightSHR(rtl)
    GENERIC MAP (178, NumberOfBits)
    PORT MAP (clk, rst, Multiplier42Weight, mbRightSHR42_Input1_56Output);

    MB_D_FF_Float_42_56_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR42_Input1_56Output, Multiplier42WeightOutput);

    InputIEEE_Float_42_56: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier42WeightOutput, flopocoMultiplier42WeightOutput);

    MB_D_FF_Float_42_56_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier42WeightOutput, flopocoMultiplier42WeightInput);

    Multiplier_Float_42: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier42WeightInput, mb_D_FF42_56MultiplierStage2Output, Multiplier42_Output_56);

    MBRightSHR_Float_42_Input2_56: entity work.MBRightSHR(rtl)
    GENERIC MAP (178, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR42_Input2_56Input, mbRightSHR42_Input2_56Output);

    MB_D_FF_Float_42_56_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR42_Input2_56Output, mb_D_FF42_56MultiplierStage1Output);

    MB_D_FF_Float_42_56_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF42_56MultiplierStage1Output, mb_D_FF42_56MultiplierStage2Output);

    MB_D_FF_Float_Adder7_Input1_14_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier42_Output_56, mb_D_FFAdder7_Input1_14_0Output);

    MB_D_FF_Float_14_57_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder7_Input1_14_0Output, mb_D_FF14_57AugendStage1Output);

    MB_D_FF_Float_14_57_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF14_57AugendStage1Output, mb_D_FF14_57AugendStage2Output);

    Adder_Float_14: entity work.FPAdd_7_24_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF14_57AugendStage2Output, mb_D_FF14_57AddendStage2Output, Adder14_Output_57);

    MB_D_FF_Float_Adder7_Input2_14_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier41_Output_55, mb_D_FFAdder7_Input2_14_0Output);

    MB_D_FF_Float_14_57_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder7_Input2_14_0Output, mb_D_FF14_57AddendStage1Output);

    MB_D_FF_Float_14_57_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF14_57AddendStage1Output, mb_D_FF14_57AddendStage2Output);

    MB_D_FF_Float_Multiplier6_Input1_43_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder14_Output_57, mb_D_FFMultiplier6_Input1_43_0Output);

    MB_D_FF_Float_43_58_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier6_Input1_43_0Output, mb_D_FF43_58MultiplicandStage1Output);

    MB_D_FF_Float_43_58_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF43_58MultiplicandStage1Output, mb_D_FF43_58MultiplicandStage2Output);

    Multiplier_Float_43: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF43_58MultiplicandStage2Output, mb_D_FF43_58MultiplierStage2Output, Multiplier43_Output_58);

    MB_D_FF_Float_Multiplier6_Input2_43_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier40_Output_54, mb_D_FFMultiplier6_Input2_43_0Output);

    MB_D_FF_Float_43_58_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier6_Input2_43_0Output, mb_D_FF43_58MultiplierStage1Output);

    MB_D_FF_Float_43_58_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF43_58MultiplierStage1Output, mb_D_FF43_58MultiplierStage2Output);

    MBRightSHR_Float_44_Input159: entity work.MBRightSHR(rtl)
    GENERIC MAP (190, NumberOfBits)
    PORT MAP (clk, rst, Multiplier44Weight, mbRightSHR44_Input1_59Output);

    MB_D_FF_Float_44_59_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR44_Input1_59Output, Multiplier44WeightOutput);

    InputIEEE_Float_44_59: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier44WeightOutput, flopocoMultiplier44WeightOutput);

    MB_D_FF_Float_44_59_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier44WeightOutput, flopocoMultiplier44WeightInput);

    Multiplier_Float_44: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier44WeightInput, mb_D_FF44_59MultiplierStage2Output, Multiplier44_Output_59);

    MBRightSHR_Float_44_Input2_59: entity work.MBRightSHR(rtl)
    GENERIC MAP (190, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR44_Input2_59Input, mbRightSHR44_Input2_59Output);

    MB_D_FF_Float_44_59_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR44_Input2_59Output, mb_D_FF44_59MultiplierStage1Output);

    MB_D_FF_Float_44_59_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF44_59MultiplierStage1Output, mb_D_FF44_59MultiplierStage2Output);

    MBRightSHR_Float_45_Input160: entity work.MBRightSHR(rtl)
    GENERIC MAP (190, NumberOfBits)
    PORT MAP (clk, rst, Multiplier45Weight, mbRightSHR45_Input1_60Output);

    MB_D_FF_Float_45_60_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR45_Input1_60Output, Multiplier45WeightOutput);

    InputIEEE_Float_45_60: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier45WeightOutput, flopocoMultiplier45WeightOutput);

    MB_D_FF_Float_45_60_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier45WeightOutput, flopocoMultiplier45WeightInput);

    Multiplier_Float_45: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier45WeightInput, mb_D_FF45_60MultiplierStage2Output, Multiplier45_Output_60);

    MBRightSHR_Float_45_Input2_60: entity work.MBRightSHR(rtl)
    GENERIC MAP (190, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR45_Input2_60Input, mbRightSHR45_Input2_60Output);

    MB_D_FF_Float_45_60_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR45_Input2_60Output, mb_D_FF45_60MultiplierStage1Output);

    MB_D_FF_Float_45_60_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF45_60MultiplierStage1Output, mb_D_FF45_60MultiplierStage2Output);

    MB_D_FF_Float_Adder6_Input1_15_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier45_Output_60, mb_D_FFAdder6_Input1_15_0Output);

    MB_D_FF_Float_15_61_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder6_Input1_15_0Output, mb_D_FF15_61AugendStage1Output);

    MB_D_FF_Float_15_61_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF15_61AugendStage1Output, mb_D_FF15_61AugendStage2Output);

    Adder_Float_15: entity work.FPAdd_7_24_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF15_61AugendStage2Output, mb_D_FF15_61AddendStage2Output, Adder15_Output_61);

    MB_D_FF_Float_Adder6_Input2_15_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier44_Output_59, mb_D_FFAdder6_Input2_15_0Output);

    MB_D_FF_Float_15_61_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder6_Input2_15_0Output, mb_D_FF15_61AddendStage1Output);

    MB_D_FF_Float_15_61_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF15_61AddendStage1Output, mb_D_FF15_61AddendStage2Output);

    MB_D_FF_Float_Multiplier5_Input1_46_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder15_Output_61, mb_D_FFMultiplier5_Input1_46_0Output);

    MB_D_FF_Float_46_62_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier5_Input1_46_0Output, mb_D_FF46_62MultiplicandStage1Output);

    MB_D_FF_Float_46_62_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF46_62MultiplicandStage1Output, mb_D_FF46_62MultiplicandStage2Output);

    Multiplier_Float_46: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF46_62MultiplicandStage2Output, mb_D_FF46_62MultiplierStage2Output, Multiplier46_Output_62);

    MB_D_FF_Float_Multiplier5_Input2_46_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier43_Output_58, mb_D_FFMultiplier5_Input2_46_0Output);

    MB_D_FF_Float_46_62_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier5_Input2_46_0Output, mb_D_FF46_62MultiplierStage1Output);

    MB_D_FF_Float_46_62_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF46_62MultiplierStage1Output, mb_D_FF46_62MultiplierStage2Output);

    MBRightSHR_Float_47_Input163: entity work.MBRightSHR(rtl)
    GENERIC MAP (202, NumberOfBits)
    PORT MAP (clk, rst, Multiplier47Weight, mbRightSHR47_Input1_63Output);

    MB_D_FF_Float_47_63_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR47_Input1_63Output, Multiplier47WeightOutput);

    InputIEEE_Float_47_63: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier47WeightOutput, flopocoMultiplier47WeightOutput);

    MB_D_FF_Float_47_63_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier47WeightOutput, flopocoMultiplier47WeightInput);

    Multiplier_Float_47: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier47WeightInput, mb_D_FF47_63MultiplierStage2Output, Multiplier47_Output_63);

    MBRightSHR_Float_47_Input2_63: entity work.MBRightSHR(rtl)
    GENERIC MAP (202, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR47_Input2_63Input, mbRightSHR47_Input2_63Output);

    MB_D_FF_Float_47_63_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR47_Input2_63Output, mb_D_FF47_63MultiplierStage1Output);

    MB_D_FF_Float_47_63_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF47_63MultiplierStage1Output, mb_D_FF47_63MultiplierStage2Output);

    MBRightSHR_Float_48_Input164: entity work.MBRightSHR(rtl)
    GENERIC MAP (202, NumberOfBits)
    PORT MAP (clk, rst, Multiplier48Weight, mbRightSHR48_Input1_64Output);

    MB_D_FF_Float_48_64_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR48_Input1_64Output, Multiplier48WeightOutput);

    InputIEEE_Float_48_64: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier48WeightOutput, flopocoMultiplier48WeightOutput);

    MB_D_FF_Float_48_64_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier48WeightOutput, flopocoMultiplier48WeightInput);

    Multiplier_Float_48: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier48WeightInput, mb_D_FF48_64MultiplierStage2Output, Multiplier48_Output_64);

    MBRightSHR_Float_48_Input2_64: entity work.MBRightSHR(rtl)
    GENERIC MAP (202, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR48_Input2_64Input, mbRightSHR48_Input2_64Output);

    MB_D_FF_Float_48_64_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR48_Input2_64Output, mb_D_FF48_64MultiplierStage1Output);

    MB_D_FF_Float_48_64_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF48_64MultiplierStage1Output, mb_D_FF48_64MultiplierStage2Output);

    MB_D_FF_Float_Adder5_Input1_16_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier48_Output_64, mb_D_FFAdder5_Input1_16_0Output);

    MB_D_FF_Float_16_65_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder5_Input1_16_0Output, mb_D_FF16_65AugendStage1Output);

    MB_D_FF_Float_16_65_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF16_65AugendStage1Output, mb_D_FF16_65AugendStage2Output);

    Adder_Float_16: entity work.FPAdd_7_24_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF16_65AugendStage2Output, mb_D_FF16_65AddendStage2Output, Adder16_Output_65);

    MB_D_FF_Float_Adder5_Input2_16_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier47_Output_63, mb_D_FFAdder5_Input2_16_0Output);

    MB_D_FF_Float_16_65_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder5_Input2_16_0Output, mb_D_FF16_65AddendStage1Output);

    MB_D_FF_Float_16_65_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF16_65AddendStage1Output, mb_D_FF16_65AddendStage2Output);

    MB_D_FF_Float_Multiplier4_Input1_49_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder16_Output_65, mb_D_FFMultiplier4_Input1_49_0Output);

    MB_D_FF_Float_49_66_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier4_Input1_49_0Output, mb_D_FF49_66MultiplicandStage1Output);

    MB_D_FF_Float_49_66_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF49_66MultiplicandStage1Output, mb_D_FF49_66MultiplicandStage2Output);

    Multiplier_Float_49: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF49_66MultiplicandStage2Output, mb_D_FF49_66MultiplierStage2Output, Multiplier49_Output_66);

    MB_D_FF_Float_Multiplier4_Input2_49_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier46_Output_62, mb_D_FFMultiplier4_Input2_49_0Output);

    MB_D_FF_Float_49_66_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier4_Input2_49_0Output, mb_D_FF49_66MultiplierStage1Output);

    MB_D_FF_Float_49_66_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF49_66MultiplierStage1Output, mb_D_FF49_66MultiplierStage2Output);

    MBRightSHR_Float_50_Input167: entity work.MBRightSHR(rtl)
    GENERIC MAP (214, NumberOfBits)
    PORT MAP (clk, rst, Multiplier50Weight, mbRightSHR50_Input1_67Output);

    MB_D_FF_Float_50_67_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR50_Input1_67Output, Multiplier50WeightOutput);

    InputIEEE_Float_50_67: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier50WeightOutput, flopocoMultiplier50WeightOutput);

    MB_D_FF_Float_50_67_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier50WeightOutput, flopocoMultiplier50WeightInput);

    Multiplier_Float_50: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier50WeightInput, mb_D_FF50_67MultiplierStage2Output, Multiplier50_Output_67);

    MBRightSHR_Float_50_Input2_67: entity work.MBRightSHR(rtl)
    GENERIC MAP (214, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR50_Input2_67Input, mbRightSHR50_Input2_67Output);

    MB_D_FF_Float_50_67_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR50_Input2_67Output, mb_D_FF50_67MultiplierStage1Output);

    MB_D_FF_Float_50_67_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF50_67MultiplierStage1Output, mb_D_FF50_67MultiplierStage2Output);

    MBRightSHR_Float_51_Input168: entity work.MBRightSHR(rtl)
    GENERIC MAP (214, NumberOfBits)
    PORT MAP (clk, rst, Multiplier51Weight, mbRightSHR51_Input1_68Output);

    MB_D_FF_Float_51_68_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR51_Input1_68Output, Multiplier51WeightOutput);

    InputIEEE_Float_51_68: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier51WeightOutput, flopocoMultiplier51WeightOutput);

    MB_D_FF_Float_51_68_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier51WeightOutput, flopocoMultiplier51WeightInput);

    Multiplier_Float_51: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier51WeightInput, mb_D_FF51_68MultiplierStage2Output, Multiplier51_Output_68);

    MBRightSHR_Float_51_Input2_68: entity work.MBRightSHR(rtl)
    GENERIC MAP (214, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR51_Input2_68Input, mbRightSHR51_Input2_68Output);

    MB_D_FF_Float_51_68_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR51_Input2_68Output, mb_D_FF51_68MultiplierStage1Output);

    MB_D_FF_Float_51_68_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF51_68MultiplierStage1Output, mb_D_FF51_68MultiplierStage2Output);

    MB_D_FF_Float_Adder4_Input1_17_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier51_Output_68, mb_D_FFAdder4_Input1_17_0Output);

    MB_D_FF_Float_17_69_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder4_Input1_17_0Output, mb_D_FF17_69AugendStage1Output);

    MB_D_FF_Float_17_69_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF17_69AugendStage1Output, mb_D_FF17_69AugendStage2Output);

    Adder_Float_17: entity work.FPAdd_7_24_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF17_69AugendStage2Output, mb_D_FF17_69AddendStage2Output, Adder17_Output_69);

    MB_D_FF_Float_Adder4_Input2_17_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier50_Output_67, mb_D_FFAdder4_Input2_17_0Output);

    MB_D_FF_Float_17_69_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder4_Input2_17_0Output, mb_D_FF17_69AddendStage1Output);

    MB_D_FF_Float_17_69_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF17_69AddendStage1Output, mb_D_FF17_69AddendStage2Output);

    MB_D_FF_Float_Multiplier3_Input1_52_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder17_Output_69, mb_D_FFMultiplier3_Input1_52_0Output);

    MB_D_FF_Float_52_70_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier3_Input1_52_0Output, mb_D_FF52_70MultiplicandStage1Output);

    MB_D_FF_Float_52_70_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF52_70MultiplicandStage1Output, mb_D_FF52_70MultiplicandStage2Output);

    Multiplier_Float_52: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF52_70MultiplicandStage2Output, mb_D_FF52_70MultiplierStage2Output, Multiplier52_Output_70);

    MB_D_FF_Float_Multiplier3_Input2_52_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier49_Output_66, mb_D_FFMultiplier3_Input2_52_0Output);

    MB_D_FF_Float_52_70_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier3_Input2_52_0Output, mb_D_FF52_70MultiplierStage1Output);

    MB_D_FF_Float_52_70_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF52_70MultiplierStage1Output, mb_D_FF52_70MultiplierStage2Output);

    MB_D_FF_Float_Multiplier2_53_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier52_Output_70, mb_D_FFMultiplier2_53_0Output);

    MB_D_FF_Float_53_71_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier2_53_0Output, mb_D_FF53_71MultiplierStage1Output);

    MB_D_FF_Float_53_71_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF53_71MultiplierStage1Output, mb_D_FF53_71MultiplierStage2Output);

    Multiplier_Float_53: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF53_71MultiplierStage2Output, flopocoMultiplier53WeightInput, Multiplier53_Output_71);

    MBRightSHR_Float_53_71: entity work.MBRightSHR(rtl)
    GENERIC MAP (250, NumberOfBits)
    PORT MAP (clk, rst, Multiplier53Weight, mbRightSHR53_71Output);

    MB_D_FF_Float_53_71_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR53_71Output, Multiplier53WeightOutput);

    InputIEEE_Float_53_71: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier53WeightOutput, flopocoMultiplier53WeightOutput);

    MB_D_FF_Float_53_71_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier53WeightOutput, flopocoMultiplier53WeightInput);

    MBRightSHR_Float_54_72: entity work.MBRightSHR(rtl)
    GENERIC MAP (4, NumberOfBits)
    PORT MAP (clk, rst, Multiplier54Weight, mbRightSHR54_72Output);

    MB_D_FF_Float_54_72_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR54_72Output, Multiplier54WeightOutput);

    InputIEEE_Float_54_72: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier54WeightOutput, flopocoMultiplier54WeightOutput);

    MB_D_FF_Float_54_72_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier54WeightOutput, flopocoMultiplier54WeightInput);

    Multiplier_Float_54: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier54WeightInput, mb_D_FF54_72MultiplierStage2Output, Multiplier54_Output_72);

    MB_D_FF_Float_Multiplier20_54_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier20_54_0Input, mb_D_FFMultiplier20_54_0Output);

    MB_D_FF_Float_54_72_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier20_54_0Output, mb_D_FF54_72MultiplierStage1Output);

    MB_D_FF_Float_54_72_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF54_72MultiplierStage1Output, mb_D_FF54_72MultiplierStage2Output);

    MBRightSHR_Float_55_73: entity work.MBRightSHR(rtl)
    GENERIC MAP (4, NumberOfBits)
    PORT MAP (clk, rst, Multiplier55Weight, mbRightSHR55_73Output);

    MB_D_FF_Float_55_73_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR55_73Output, Multiplier55WeightOutput);

    InputIEEE_Float_55_73: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier55WeightOutput, flopocoMultiplier55WeightOutput);

    MB_D_FF_Float_55_73_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier55WeightOutput, flopocoMultiplier55WeightInput);

    Multiplier_Float_55: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier55WeightInput, mb_D_FF55_73MultiplierStage2Output, Multiplier55_Output_73);

    MB_D_FF_Float_Multiplier20_55_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier20_55_0Input, mb_D_FFMultiplier20_55_0Output);

    MB_D_FF_Float_55_73_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier20_55_0Output, mb_D_FF55_73MultiplierStage1Output);

    MB_D_FF_Float_55_73_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF55_73MultiplierStage1Output, mb_D_FF55_73MultiplierStage2Output);

    MB_D_FF_Float_Adder19_Input1_18_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier55_Output_73, mb_D_FFAdder19_Input1_18_0Output);

    MB_D_FF_Float_18_74_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder19_Input1_18_0Output, mb_D_FF18_74AugendStage1Output);

    MB_D_FF_Float_18_74_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF18_74AugendStage1Output, mb_D_FF18_74AugendStage2Output);

    Adder_Float_18: entity work.FPAdd_7_24_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF18_74AugendStage2Output, mb_D_FF18_74AddendStage2Output, Adder18_Output_74);

    MB_D_FF_Float_Adder19_Input2_18_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier54_Output_72, mb_D_FFAdder19_Input2_18_0Output);

    MB_D_FF_Float_18_74_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder19_Input2_18_0Output, mb_D_FF18_74AddendStage1Output);

    MB_D_FF_Float_18_74_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF18_74AddendStage1Output, mb_D_FF18_74AddendStage2Output);

    MBRightSHR_Float_56_75: entity work.MBRightSHR(rtl)
    GENERIC MAP (4, NumberOfBits)
    PORT MAP (clk, rst, Multiplier56Weight, mbRightSHR56_75Output);

    MB_D_FF_Float_56_75_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR56_75Output, Multiplier56WeightOutput);

    InputIEEE_Float_56_75: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier56WeightOutput, flopocoMultiplier56WeightOutput);

    MB_D_FF_Float_56_75_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier56WeightOutput, flopocoMultiplier56WeightInput);

    Multiplier_Float_56: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier56WeightInput, mb_D_FF56_75MultiplierStage2Output, Multiplier56_Output_75);

    MB_D_FF_Float_Multiplier20_56_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier20_56_0Input, mb_D_FFMultiplier20_56_0Output);

    MB_D_FF_Float_56_75_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier20_56_0Output, mb_D_FF56_75MultiplierStage1Output);

    MB_D_FF_Float_56_75_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF56_75MultiplierStage1Output, mb_D_FF56_75MultiplierStage2Output);

    MBRightSHR_Float_57_76: entity work.MBRightSHR(rtl)
    GENERIC MAP (4, NumberOfBits)
    PORT MAP (clk, rst, Multiplier57Weight, mbRightSHR57_76Output);

    MB_D_FF_Float_57_76_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR57_76Output, Multiplier57WeightOutput);

    InputIEEE_Float_57_76: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier57WeightOutput, flopocoMultiplier57WeightOutput);

    MB_D_FF_Float_57_76_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier57WeightOutput, flopocoMultiplier57WeightInput);

    Multiplier_Float_57: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier57WeightInput, mb_D_FF57_76MultiplierStage2Output, Multiplier57_Output_76);

    MB_D_FF_Float_Multiplier20_57_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier20_57_0Input, mb_D_FFMultiplier20_57_0Output);

    MB_D_FF_Float_57_76_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier20_57_0Output, mb_D_FF57_76MultiplierStage1Output);

    MB_D_FF_Float_57_76_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF57_76MultiplierStage1Output, mb_D_FF57_76MultiplierStage2Output);

    MB_D_FF_Float_Adder19_Input1_19_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier57_Output_76, mb_D_FFAdder19_Input1_19_0Output);

    MB_D_FF_Float_19_77_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder19_Input1_19_0Output, mb_D_FF19_77AugendStage1Output);

    MB_D_FF_Float_19_77_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF19_77AugendStage1Output, mb_D_FF19_77AugendStage2Output);

    Adder_Float_19: entity work.FPAdd_7_24_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF19_77AugendStage2Output, mb_D_FF19_77AddendStage2Output, Adder19_Output_77);

    MB_D_FF_Float_Adder19_Input2_19_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier56_Output_75, mb_D_FFAdder19_Input2_19_0Output);

    MB_D_FF_Float_19_77_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder19_Input2_19_0Output, mb_D_FF19_77AddendStage1Output);

    MB_D_FF_Float_19_77_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF19_77AddendStage1Output, mb_D_FF19_77AddendStage2Output);

    MB_D_FF_Float_Multiplier18_Input1_58_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder19_Output_77, mb_D_FFMultiplier18_Input1_58_0Output);

    MB_D_FF_Float_58_78_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier18_Input1_58_0Output, mb_D_FF58_78MultiplicandStage1Output);

    MB_D_FF_Float_58_78_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF58_78MultiplicandStage1Output, mb_D_FF58_78MultiplicandStage2Output);

    Multiplier_Float_58: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF58_78MultiplicandStage2Output, mb_D_FF58_78MultiplierStage2Output, Multiplier58_Output_78);

    MB_D_FF_Float_Multiplier18_Input2_58_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder18_Output_74, mb_D_FFMultiplier18_Input2_58_0Output);

    MB_D_FF_Float_58_78_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier18_Input2_58_0Output, mb_D_FF58_78MultiplierStage1Output);

    MB_D_FF_Float_58_78_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF58_78MultiplierStage1Output, mb_D_FF58_78MultiplierStage2Output);

    MBRightSHR_Float_59_Input179: entity work.MBRightSHR(rtl)
    GENERIC MAP (16, NumberOfBits)
    PORT MAP (clk, rst, Multiplier59Weight, mbRightSHR59_Input1_79Output);

    MB_D_FF_Float_59_79_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR59_Input1_79Output, Multiplier59WeightOutput);

    InputIEEE_Float_59_79: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier59WeightOutput, flopocoMultiplier59WeightOutput);

    MB_D_FF_Float_59_79_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier59WeightOutput, flopocoMultiplier59WeightInput);

    Multiplier_Float_59: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier59WeightInput, mb_D_FF59_79MultiplierStage2Output, Multiplier59_Output_79);

    MBRightSHR_Float_59_Input2_79: entity work.MBRightSHR(rtl)
    GENERIC MAP (16, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR59_Input2_79Input, mbRightSHR59_Input2_79Output);

    MB_D_FF_Float_59_79_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR59_Input2_79Output, mb_D_FF59_79MultiplierStage1Output);

    MB_D_FF_Float_59_79_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF59_79MultiplierStage1Output, mb_D_FF59_79MultiplierStage2Output);

    MBRightSHR_Float_60_Input180: entity work.MBRightSHR(rtl)
    GENERIC MAP (16, NumberOfBits)
    PORT MAP (clk, rst, Multiplier60Weight, mbRightSHR60_Input1_80Output);

    MB_D_FF_Float_60_80_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR60_Input1_80Output, Multiplier60WeightOutput);

    InputIEEE_Float_60_80: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier60WeightOutput, flopocoMultiplier60WeightOutput);

    MB_D_FF_Float_60_80_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier60WeightOutput, flopocoMultiplier60WeightInput);

    Multiplier_Float_60: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier60WeightInput, mb_D_FF60_80MultiplierStage2Output, Multiplier60_Output_80);

    MBRightSHR_Float_60_Input2_80: entity work.MBRightSHR(rtl)
    GENERIC MAP (16, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR60_Input2_80Input, mbRightSHR60_Input2_80Output);

    MB_D_FF_Float_60_80_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR60_Input2_80Output, mb_D_FF60_80MultiplierStage1Output);

    MB_D_FF_Float_60_80_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF60_80MultiplierStage1Output, mb_D_FF60_80MultiplierStage2Output);

    MB_D_FF_Float_Adder18_Input1_20_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier60_Output_80, mb_D_FFAdder18_Input1_20_0Output);

    MB_D_FF_Float_20_81_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder18_Input1_20_0Output, mb_D_FF20_81AugendStage1Output);

    MB_D_FF_Float_20_81_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF20_81AugendStage1Output, mb_D_FF20_81AugendStage2Output);

    Adder_Float_20: entity work.FPAdd_7_24_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF20_81AugendStage2Output, mb_D_FF20_81AddendStage2Output, Adder20_Output_81);

    MB_D_FF_Float_Adder18_Input2_20_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier59_Output_79, mb_D_FFAdder18_Input2_20_0Output);

    MB_D_FF_Float_20_81_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder18_Input2_20_0Output, mb_D_FF20_81AddendStage1Output);

    MB_D_FF_Float_20_81_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF20_81AddendStage1Output, mb_D_FF20_81AddendStage2Output);

    MB_D_FF_Float_Multiplier17_Input1_61_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder20_Output_81, mb_D_FFMultiplier17_Input1_61_0Output);

    MB_D_FF_Float_61_82_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier17_Input1_61_0Output, mb_D_FF61_82MultiplicandStage1Output);

    MB_D_FF_Float_61_82_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF61_82MultiplicandStage1Output, mb_D_FF61_82MultiplicandStage2Output);

    Multiplier_Float_61: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF61_82MultiplicandStage2Output, mb_D_FF61_82MultiplierStage2Output, Multiplier61_Output_82);

    MB_D_FF_Float_Multiplier17_Input2_61_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier58_Output_78, mb_D_FFMultiplier17_Input2_61_0Output);

    MB_D_FF_Float_61_82_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier17_Input2_61_0Output, mb_D_FF61_82MultiplierStage1Output);

    MB_D_FF_Float_61_82_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF61_82MultiplierStage1Output, mb_D_FF61_82MultiplierStage2Output);

    MBRightSHR_Float_62_Input183: entity work.MBRightSHR(rtl)
    GENERIC MAP (43, NumberOfBits)
    PORT MAP (clk, rst, Multiplier62Weight, mbRightSHR62_Input1_83Output);

    MB_D_FF_Float_62_83_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR62_Input1_83Output, Multiplier62WeightOutput);

    InputIEEE_Float_62_83: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier62WeightOutput, flopocoMultiplier62WeightOutput);

    MB_D_FF_Float_62_83_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier62WeightOutput, flopocoMultiplier62WeightInput);

    Multiplier_Float_62: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier62WeightInput, mb_D_FF62_83MultiplierStage2Output, Multiplier62_Output_83);

    MBRightSHR_Float_62_Input2_83: entity work.MBRightSHR(rtl)
    GENERIC MAP (43, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR62_Input2_83Input, mbRightSHR62_Input2_83Output);

    MB_D_FF_Float_62_83_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR62_Input2_83Output, mb_D_FF62_83MultiplierStage1Output);

    MB_D_FF_Float_62_83_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF62_83MultiplierStage1Output, mb_D_FF62_83MultiplierStage2Output);

    MBRightSHR_Float_63_Input184: entity work.MBRightSHR(rtl)
    GENERIC MAP (43, NumberOfBits)
    PORT MAP (clk, rst, Multiplier63Weight, mbRightSHR63_Input1_84Output);

    MB_D_FF_Float_63_84_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR63_Input1_84Output, Multiplier63WeightOutput);

    InputIEEE_Float_63_84: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier63WeightOutput, flopocoMultiplier63WeightOutput);

    MB_D_FF_Float_63_84_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier63WeightOutput, flopocoMultiplier63WeightInput);

    Multiplier_Float_63: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier63WeightInput, mb_D_FF63_84MultiplierStage2Output, Multiplier63_Output_84);

    MBRightSHR_Float_63_Input2_84: entity work.MBRightSHR(rtl)
    GENERIC MAP (43, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR63_Input2_84Input, mbRightSHR63_Input2_84Output);

    MB_D_FF_Float_63_84_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR63_Input2_84Output, mb_D_FF63_84MultiplierStage1Output);

    MB_D_FF_Float_63_84_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF63_84MultiplierStage1Output, mb_D_FF63_84MultiplierStage2Output);

    MB_D_FF_Float_Adder17_Input1_21_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier63_Output_84, mb_D_FFAdder17_Input1_21_0Output);

    MB_D_FF_Float_21_85_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder17_Input1_21_0Output, mb_D_FF21_85AugendStage1Output);

    MB_D_FF_Float_21_85_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF21_85AugendStage1Output, mb_D_FF21_85AugendStage2Output);

    Adder_Float_21: entity work.FPAdd_7_24_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF21_85AugendStage2Output, mb_D_FF21_85AddendStage2Output, Adder21_Output_85);

    MB_D_FF_Float_Adder17_Input2_21_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier62_Output_83, mb_D_FFAdder17_Input2_21_0Output);

    MB_D_FF_Float_21_85_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder17_Input2_21_0Output, mb_D_FF21_85AddendStage1Output);

    MB_D_FF_Float_21_85_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF21_85AddendStage1Output, mb_D_FF21_85AddendStage2Output);

    MB_D_FF_Float_Multiplier16_Input1_64_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder21_Output_85, mb_D_FFMultiplier16_Input1_64_0Output);

    MB_D_FF_Float_64_86_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier16_Input1_64_0Output, mb_D_FF64_86MultiplicandStage1Output);

    MB_D_FF_Float_64_86_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF64_86MultiplicandStage1Output, mb_D_FF64_86MultiplicandStage2Output);

    Multiplier_Float_64: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF64_86MultiplicandStage2Output, mb_D_FF64_86MultiplierStage2Output, Multiplier64_Output_86);

    MB_D_FF_Float_Multiplier16_Input2_64_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier61_Output_82, mb_D_FFMultiplier16_Input2_64_0Output);

    MB_D_FF_Float_64_86_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier16_Input2_64_0Output, mb_D_FF64_86MultiplierStage1Output);

    MB_D_FF_Float_64_86_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF64_86MultiplierStage1Output, mb_D_FF64_86MultiplierStage2Output);

    MBRightSHR_Float_65_Input187: entity work.MBRightSHR(rtl)
    GENERIC MAP (55, NumberOfBits)
    PORT MAP (clk, rst, Multiplier65Weight, mbRightSHR65_Input1_87Output);

    MB_D_FF_Float_65_87_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR65_Input1_87Output, Multiplier65WeightOutput);

    InputIEEE_Float_65_87: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier65WeightOutput, flopocoMultiplier65WeightOutput);

    MB_D_FF_Float_65_87_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier65WeightOutput, flopocoMultiplier65WeightInput);

    Multiplier_Float_65: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier65WeightInput, mb_D_FF65_87MultiplierStage2Output, Multiplier65_Output_87);

    MBRightSHR_Float_65_Input2_87: entity work.MBRightSHR(rtl)
    GENERIC MAP (55, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR65_Input2_87Input, mbRightSHR65_Input2_87Output);

    MB_D_FF_Float_65_87_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR65_Input2_87Output, mb_D_FF65_87MultiplierStage1Output);

    MB_D_FF_Float_65_87_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF65_87MultiplierStage1Output, mb_D_FF65_87MultiplierStage2Output);

    MBRightSHR_Float_66_Input188: entity work.MBRightSHR(rtl)
    GENERIC MAP (55, NumberOfBits)
    PORT MAP (clk, rst, Multiplier66Weight, mbRightSHR66_Input1_88Output);

    MB_D_FF_Float_66_88_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR66_Input1_88Output, Multiplier66WeightOutput);

    InputIEEE_Float_66_88: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier66WeightOutput, flopocoMultiplier66WeightOutput);

    MB_D_FF_Float_66_88_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier66WeightOutput, flopocoMultiplier66WeightInput);

    Multiplier_Float_66: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier66WeightInput, mb_D_FF66_88MultiplierStage2Output, Multiplier66_Output_88);

    MBRightSHR_Float_66_Input2_88: entity work.MBRightSHR(rtl)
    GENERIC MAP (55, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR66_Input2_88Input, mbRightSHR66_Input2_88Output);

    MB_D_FF_Float_66_88_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR66_Input2_88Output, mb_D_FF66_88MultiplierStage1Output);

    MB_D_FF_Float_66_88_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF66_88MultiplierStage1Output, mb_D_FF66_88MultiplierStage2Output);

    MB_D_FF_Float_Adder16_Input1_22_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier66_Output_88, mb_D_FFAdder16_Input1_22_0Output);

    MB_D_FF_Float_22_89_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder16_Input1_22_0Output, mb_D_FF22_89AugendStage1Output);

    MB_D_FF_Float_22_89_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF22_89AugendStage1Output, mb_D_FF22_89AugendStage2Output);

    Adder_Float_22: entity work.FPAdd_7_24_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF22_89AugendStage2Output, mb_D_FF22_89AddendStage2Output, Adder22_Output_89);

    MB_D_FF_Float_Adder16_Input2_22_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier65_Output_87, mb_D_FFAdder16_Input2_22_0Output);

    MB_D_FF_Float_22_89_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder16_Input2_22_0Output, mb_D_FF22_89AddendStage1Output);

    MB_D_FF_Float_22_89_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF22_89AddendStage1Output, mb_D_FF22_89AddendStage2Output);

    MB_D_FF_Float_Multiplier15_Input1_67_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder22_Output_89, mb_D_FFMultiplier15_Input1_67_0Output);

    MB_D_FF_Float_67_90_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier15_Input1_67_0Output, mb_D_FF67_90MultiplicandStage1Output);

    MB_D_FF_Float_67_90_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF67_90MultiplicandStage1Output, mb_D_FF67_90MultiplicandStage2Output);

    Multiplier_Float_67: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF67_90MultiplicandStage2Output, mb_D_FF67_90MultiplierStage2Output, Multiplier67_Output_90);

    MB_D_FF_Float_Multiplier15_Input2_67_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier64_Output_86, mb_D_FFMultiplier15_Input2_67_0Output);

    MB_D_FF_Float_67_90_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier15_Input2_67_0Output, mb_D_FF67_90MultiplierStage1Output);

    MB_D_FF_Float_67_90_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF67_90MultiplierStage1Output, mb_D_FF67_90MultiplierStage2Output);

    MBRightSHR_Float_68_Input191: entity work.MBRightSHR(rtl)
    GENERIC MAP (67, NumberOfBits)
    PORT MAP (clk, rst, Multiplier68Weight, mbRightSHR68_Input1_91Output);

    MB_D_FF_Float_68_91_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR68_Input1_91Output, Multiplier68WeightOutput);

    InputIEEE_Float_68_91: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier68WeightOutput, flopocoMultiplier68WeightOutput);

    MB_D_FF_Float_68_91_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier68WeightOutput, flopocoMultiplier68WeightInput);

    Multiplier_Float_68: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier68WeightInput, mb_D_FF68_91MultiplierStage2Output, Multiplier68_Output_91);

    MBRightSHR_Float_68_Input2_91: entity work.MBRightSHR(rtl)
    GENERIC MAP (67, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR68_Input2_91Input, mbRightSHR68_Input2_91Output);

    MB_D_FF_Float_68_91_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR68_Input2_91Output, mb_D_FF68_91MultiplierStage1Output);

    MB_D_FF_Float_68_91_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF68_91MultiplierStage1Output, mb_D_FF68_91MultiplierStage2Output);

    MBRightSHR_Float_69_Input192: entity work.MBRightSHR(rtl)
    GENERIC MAP (67, NumberOfBits)
    PORT MAP (clk, rst, Multiplier69Weight, mbRightSHR69_Input1_92Output);

    MB_D_FF_Float_69_92_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR69_Input1_92Output, Multiplier69WeightOutput);

    InputIEEE_Float_69_92: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier69WeightOutput, flopocoMultiplier69WeightOutput);

    MB_D_FF_Float_69_92_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier69WeightOutput, flopocoMultiplier69WeightInput);

    Multiplier_Float_69: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier69WeightInput, mb_D_FF69_92MultiplierStage2Output, Multiplier69_Output_92);

    MBRightSHR_Float_69_Input2_92: entity work.MBRightSHR(rtl)
    GENERIC MAP (67, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR69_Input2_92Input, mbRightSHR69_Input2_92Output);

    MB_D_FF_Float_69_92_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR69_Input2_92Output, mb_D_FF69_92MultiplierStage1Output);

    MB_D_FF_Float_69_92_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF69_92MultiplierStage1Output, mb_D_FF69_92MultiplierStage2Output);

    MB_D_FF_Float_Adder15_Input1_23_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier69_Output_92, mb_D_FFAdder15_Input1_23_0Output);

    MB_D_FF_Float_23_93_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder15_Input1_23_0Output, mb_D_FF23_93AugendStage1Output);

    MB_D_FF_Float_23_93_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF23_93AugendStage1Output, mb_D_FF23_93AugendStage2Output);

    Adder_Float_23: entity work.FPAdd_7_24_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF23_93AugendStage2Output, mb_D_FF23_93AddendStage2Output, Adder23_Output_93);

    MB_D_FF_Float_Adder15_Input2_23_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier68_Output_91, mb_D_FFAdder15_Input2_23_0Output);

    MB_D_FF_Float_23_93_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder15_Input2_23_0Output, mb_D_FF23_93AddendStage1Output);

    MB_D_FF_Float_23_93_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF23_93AddendStage1Output, mb_D_FF23_93AddendStage2Output);

    MB_D_FF_Float_Multiplier14_Input1_70_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder23_Output_93, mb_D_FFMultiplier14_Input1_70_0Output);

    MB_D_FF_Float_70_94_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier14_Input1_70_0Output, mb_D_FF70_94MultiplicandStage1Output);

    MB_D_FF_Float_70_94_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF70_94MultiplicandStage1Output, mb_D_FF70_94MultiplicandStage2Output);

    Multiplier_Float_70: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF70_94MultiplicandStage2Output, mb_D_FF70_94MultiplierStage2Output, Multiplier70_Output_94);

    MB_D_FF_Float_Multiplier14_Input2_70_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier67_Output_90, mb_D_FFMultiplier14_Input2_70_0Output);

    MB_D_FF_Float_70_94_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier14_Input2_70_0Output, mb_D_FF70_94MultiplierStage1Output);

    MB_D_FF_Float_70_94_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF70_94MultiplierStage1Output, mb_D_FF70_94MultiplierStage2Output);

    MBRightSHR_Float_71_Input195: entity work.MBRightSHR(rtl)
    GENERIC MAP (94, NumberOfBits)
    PORT MAP (clk, rst, Multiplier71Weight, mbRightSHR71_Input1_95Output);

    MB_D_FF_Float_71_95_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR71_Input1_95Output, Multiplier71WeightOutput);

    InputIEEE_Float_71_95: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier71WeightOutput, flopocoMultiplier71WeightOutput);

    MB_D_FF_Float_71_95_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier71WeightOutput, flopocoMultiplier71WeightInput);

    Multiplier_Float_71: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier71WeightInput, mb_D_FF71_95MultiplierStage2Output, Multiplier71_Output_95);

    MBRightSHR_Float_71_Input2_95: entity work.MBRightSHR(rtl)
    GENERIC MAP (94, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR71_Input2_95Input, mbRightSHR71_Input2_95Output);

    MB_D_FF_Float_71_95_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR71_Input2_95Output, mb_D_FF71_95MultiplierStage1Output);

    MB_D_FF_Float_71_95_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF71_95MultiplierStage1Output, mb_D_FF71_95MultiplierStage2Output);

    MBRightSHR_Float_72_Input196: entity work.MBRightSHR(rtl)
    GENERIC MAP (94, NumberOfBits)
    PORT MAP (clk, rst, Multiplier72Weight, mbRightSHR72_Input1_96Output);

    MB_D_FF_Float_72_96_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR72_Input1_96Output, Multiplier72WeightOutput);

    InputIEEE_Float_72_96: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier72WeightOutput, flopocoMultiplier72WeightOutput);

    MB_D_FF_Float_72_96_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier72WeightOutput, flopocoMultiplier72WeightInput);

    Multiplier_Float_72: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier72WeightInput, mb_D_FF72_96MultiplierStage2Output, Multiplier72_Output_96);

    MBRightSHR_Float_72_Input2_96: entity work.MBRightSHR(rtl)
    GENERIC MAP (94, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR72_Input2_96Input, mbRightSHR72_Input2_96Output);

    MB_D_FF_Float_72_96_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR72_Input2_96Output, mb_D_FF72_96MultiplierStage1Output);

    MB_D_FF_Float_72_96_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF72_96MultiplierStage1Output, mb_D_FF72_96MultiplierStage2Output);

    MB_D_FF_Float_Adder14_Input1_24_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier72_Output_96, mb_D_FFAdder14_Input1_24_0Output);

    MB_D_FF_Float_24_97_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder14_Input1_24_0Output, mb_D_FF24_97AugendStage1Output);

    MB_D_FF_Float_24_97_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF24_97AugendStage1Output, mb_D_FF24_97AugendStage2Output);

    Adder_Float_24: entity work.FPAdd_7_24_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF24_97AugendStage2Output, mb_D_FF24_97AddendStage2Output, Adder24_Output_97);

    MB_D_FF_Float_Adder14_Input2_24_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier71_Output_95, mb_D_FFAdder14_Input2_24_0Output);

    MB_D_FF_Float_24_97_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder14_Input2_24_0Output, mb_D_FF24_97AddendStage1Output);

    MB_D_FF_Float_24_97_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF24_97AddendStage1Output, mb_D_FF24_97AddendStage2Output);

    MB_D_FF_Float_Multiplier13_Input1_73_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder24_Output_97, mb_D_FFMultiplier13_Input1_73_0Output);

    MB_D_FF_Float_73_98_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier13_Input1_73_0Output, mb_D_FF73_98MultiplicandStage1Output);

    MB_D_FF_Float_73_98_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF73_98MultiplicandStage1Output, mb_D_FF73_98MultiplicandStage2Output);

    Multiplier_Float_73: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF73_98MultiplicandStage2Output, mb_D_FF73_98MultiplierStage2Output, Multiplier73_Output_98);

    MB_D_FF_Float_Multiplier13_Input2_73_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier70_Output_94, mb_D_FFMultiplier13_Input2_73_0Output);

    MB_D_FF_Float_73_98_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier13_Input2_73_0Output, mb_D_FF73_98MultiplierStage1Output);

    MB_D_FF_Float_73_98_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF73_98MultiplierStage1Output, mb_D_FF73_98MultiplierStage2Output);

    MBRightSHR_Float_74_Input199: entity work.MBRightSHR(rtl)
    GENERIC MAP (106, NumberOfBits)
    PORT MAP (clk, rst, Multiplier74Weight, mbRightSHR74_Input1_99Output);

    MB_D_FF_Float_74_99_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR74_Input1_99Output, Multiplier74WeightOutput);

    InputIEEE_Float_74_99: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier74WeightOutput, flopocoMultiplier74WeightOutput);

    MB_D_FF_Float_74_99_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier74WeightOutput, flopocoMultiplier74WeightInput);

    Multiplier_Float_74: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier74WeightInput, mb_D_FF74_99MultiplierStage2Output, Multiplier74_Output_99);

    MBRightSHR_Float_74_Input2_99: entity work.MBRightSHR(rtl)
    GENERIC MAP (106, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR74_Input2_99Input, mbRightSHR74_Input2_99Output);

    MB_D_FF_Float_74_99_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR74_Input2_99Output, mb_D_FF74_99MultiplierStage1Output);

    MB_D_FF_Float_74_99_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF74_99MultiplierStage1Output, mb_D_FF74_99MultiplierStage2Output);

    MBRightSHR_Float_75_Input1100: entity work.MBRightSHR(rtl)
    GENERIC MAP (106, NumberOfBits)
    PORT MAP (clk, rst, Multiplier75Weight, mbRightSHR75_Input1_100Output);

    MB_D_FF_Float_75_100_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR75_Input1_100Output, Multiplier75WeightOutput);

    InputIEEE_Float_75_100: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier75WeightOutput, flopocoMultiplier75WeightOutput);

    MB_D_FF_Float_75_100_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier75WeightOutput, flopocoMultiplier75WeightInput);

    Multiplier_Float_75: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier75WeightInput, mb_D_FF75_100MultiplierStage2Output, Multiplier75_Output_100);

    MBRightSHR_Float_75_Input2_100: entity work.MBRightSHR(rtl)
    GENERIC MAP (106, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR75_Input2_100Input, mbRightSHR75_Input2_100Output);

    MB_D_FF_Float_75_100_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR75_Input2_100Output, mb_D_FF75_100MultiplierStage1Output);

    MB_D_FF_Float_75_100_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF75_100MultiplierStage1Output, mb_D_FF75_100MultiplierStage2Output);

    MB_D_FF_Float_Adder13_Input1_25_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier75_Output_100, mb_D_FFAdder13_Input1_25_0Output);

    MB_D_FF_Float_25_101_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder13_Input1_25_0Output, mb_D_FF25_101AugendStage1Output);

    MB_D_FF_Float_25_101_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF25_101AugendStage1Output, mb_D_FF25_101AugendStage2Output);

    Adder_Float_25: entity work.FPAdd_7_24_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF25_101AugendStage2Output, mb_D_FF25_101AddendStage2Output, Adder25_Output_101);

    MB_D_FF_Float_Adder13_Input2_25_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier74_Output_99, mb_D_FFAdder13_Input2_25_0Output);

    MB_D_FF_Float_25_101_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder13_Input2_25_0Output, mb_D_FF25_101AddendStage1Output);

    MB_D_FF_Float_25_101_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF25_101AddendStage1Output, mb_D_FF25_101AddendStage2Output);

    MB_D_FF_Float_Multiplier12_Input1_76_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder25_Output_101, mb_D_FFMultiplier12_Input1_76_0Output);

    MB_D_FF_Float_76_102_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier12_Input1_76_0Output, mb_D_FF76_102MultiplicandStage1Output);

    MB_D_FF_Float_76_102_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF76_102MultiplicandStage1Output, mb_D_FF76_102MultiplicandStage2Output);

    Multiplier_Float_76: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF76_102MultiplicandStage2Output, mb_D_FF76_102MultiplierStage2Output, Multiplier76_Output_102);

    MB_D_FF_Float_Multiplier12_Input2_76_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier73_Output_98, mb_D_FFMultiplier12_Input2_76_0Output);

    MB_D_FF_Float_76_102_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier12_Input2_76_0Output, mb_D_FF76_102MultiplierStage1Output);

    MB_D_FF_Float_76_102_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF76_102MultiplierStage1Output, mb_D_FF76_102MultiplierStage2Output);

    MBRightSHR_Float_77_Input1103: entity work.MBRightSHR(rtl)
    GENERIC MAP (118, NumberOfBits)
    PORT MAP (clk, rst, Multiplier77Weight, mbRightSHR77_Input1_103Output);

    MB_D_FF_Float_77_103_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR77_Input1_103Output, Multiplier77WeightOutput);

    InputIEEE_Float_77_103: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier77WeightOutput, flopocoMultiplier77WeightOutput);

    MB_D_FF_Float_77_103_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier77WeightOutput, flopocoMultiplier77WeightInput);

    Multiplier_Float_77: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier77WeightInput, mb_D_FF77_103MultiplierStage2Output, Multiplier77_Output_103);

    MBRightSHR_Float_77_Input2_103: entity work.MBRightSHR(rtl)
    GENERIC MAP (118, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR77_Input2_103Input, mbRightSHR77_Input2_103Output);

    MB_D_FF_Float_77_103_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR77_Input2_103Output, mb_D_FF77_103MultiplierStage1Output);

    MB_D_FF_Float_77_103_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF77_103MultiplierStage1Output, mb_D_FF77_103MultiplierStage2Output);

    MBRightSHR_Float_78_Input1104: entity work.MBRightSHR(rtl)
    GENERIC MAP (118, NumberOfBits)
    PORT MAP (clk, rst, Multiplier78Weight, mbRightSHR78_Input1_104Output);

    MB_D_FF_Float_78_104_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR78_Input1_104Output, Multiplier78WeightOutput);

    InputIEEE_Float_78_104: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier78WeightOutput, flopocoMultiplier78WeightOutput);

    MB_D_FF_Float_78_104_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier78WeightOutput, flopocoMultiplier78WeightInput);

    Multiplier_Float_78: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier78WeightInput, mb_D_FF78_104MultiplierStage2Output, Multiplier78_Output_104);

    MBRightSHR_Float_78_Input2_104: entity work.MBRightSHR(rtl)
    GENERIC MAP (118, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR78_Input2_104Input, mbRightSHR78_Input2_104Output);

    MB_D_FF_Float_78_104_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR78_Input2_104Output, mb_D_FF78_104MultiplierStage1Output);

    MB_D_FF_Float_78_104_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF78_104MultiplierStage1Output, mb_D_FF78_104MultiplierStage2Output);

    MB_D_FF_Float_Adder12_Input1_26_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier78_Output_104, mb_D_FFAdder12_Input1_26_0Output);

    MB_D_FF_Float_26_105_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder12_Input1_26_0Output, mb_D_FF26_105AugendStage1Output);

    MB_D_FF_Float_26_105_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF26_105AugendStage1Output, mb_D_FF26_105AugendStage2Output);

    Adder_Float_26: entity work.FPAdd_7_24_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF26_105AugendStage2Output, mb_D_FF26_105AddendStage2Output, Adder26_Output_105);

    MB_D_FF_Float_Adder12_Input2_26_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier77_Output_103, mb_D_FFAdder12_Input2_26_0Output);

    MB_D_FF_Float_26_105_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder12_Input2_26_0Output, mb_D_FF26_105AddendStage1Output);

    MB_D_FF_Float_26_105_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF26_105AddendStage1Output, mb_D_FF26_105AddendStage2Output);

    MB_D_FF_Float_Multiplier11_Input1_79_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder26_Output_105, mb_D_FFMultiplier11_Input1_79_0Output);

    MB_D_FF_Float_79_106_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier11_Input1_79_0Output, mb_D_FF79_106MultiplicandStage1Output);

    MB_D_FF_Float_79_106_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF79_106MultiplicandStage1Output, mb_D_FF79_106MultiplicandStage2Output);

    Multiplier_Float_79: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF79_106MultiplicandStage2Output, mb_D_FF79_106MultiplierStage2Output, Multiplier79_Output_106);

    MB_D_FF_Float_Multiplier11_Input2_79_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier76_Output_102, mb_D_FFMultiplier11_Input2_79_0Output);

    MB_D_FF_Float_79_106_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier11_Input2_79_0Output, mb_D_FF79_106MultiplierStage1Output);

    MB_D_FF_Float_79_106_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF79_106MultiplierStage1Output, mb_D_FF79_106MultiplierStage2Output);

    MBRightSHR_Float_80_Input1107: entity work.MBRightSHR(rtl)
    GENERIC MAP (130, NumberOfBits)
    PORT MAP (clk, rst, Multiplier80Weight, mbRightSHR80_Input1_107Output);

    MB_D_FF_Float_80_107_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR80_Input1_107Output, Multiplier80WeightOutput);

    InputIEEE_Float_80_107: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier80WeightOutput, flopocoMultiplier80WeightOutput);

    MB_D_FF_Float_80_107_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier80WeightOutput, flopocoMultiplier80WeightInput);

    Multiplier_Float_80: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier80WeightInput, mb_D_FF80_107MultiplierStage2Output, Multiplier80_Output_107);

    MBRightSHR_Float_80_Input2_107: entity work.MBRightSHR(rtl)
    GENERIC MAP (130, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR80_Input2_107Input, mbRightSHR80_Input2_107Output);

    MB_D_FF_Float_80_107_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR80_Input2_107Output, mb_D_FF80_107MultiplierStage1Output);

    MB_D_FF_Float_80_107_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF80_107MultiplierStage1Output, mb_D_FF80_107MultiplierStage2Output);

    MBRightSHR_Float_81_Input1108: entity work.MBRightSHR(rtl)
    GENERIC MAP (130, NumberOfBits)
    PORT MAP (clk, rst, Multiplier81Weight, mbRightSHR81_Input1_108Output);

    MB_D_FF_Float_81_108_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR81_Input1_108Output, Multiplier81WeightOutput);

    InputIEEE_Float_81_108: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier81WeightOutput, flopocoMultiplier81WeightOutput);

    MB_D_FF_Float_81_108_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier81WeightOutput, flopocoMultiplier81WeightInput);

    Multiplier_Float_81: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier81WeightInput, mb_D_FF81_108MultiplierStage2Output, Multiplier81_Output_108);

    MBRightSHR_Float_81_Input2_108: entity work.MBRightSHR(rtl)
    GENERIC MAP (130, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR81_Input2_108Input, mbRightSHR81_Input2_108Output);

    MB_D_FF_Float_81_108_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR81_Input2_108Output, mb_D_FF81_108MultiplierStage1Output);

    MB_D_FF_Float_81_108_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF81_108MultiplierStage1Output, mb_D_FF81_108MultiplierStage2Output);

    MB_D_FF_Float_Adder11_Input1_27_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier81_Output_108, mb_D_FFAdder11_Input1_27_0Output);

    MB_D_FF_Float_27_109_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder11_Input1_27_0Output, mb_D_FF27_109AugendStage1Output);

    MB_D_FF_Float_27_109_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF27_109AugendStage1Output, mb_D_FF27_109AugendStage2Output);

    Adder_Float_27: entity work.FPAdd_7_24_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF27_109AugendStage2Output, mb_D_FF27_109AddendStage2Output, Adder27_Output_109);

    MB_D_FF_Float_Adder11_Input2_27_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier80_Output_107, mb_D_FFAdder11_Input2_27_0Output);

    MB_D_FF_Float_27_109_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder11_Input2_27_0Output, mb_D_FF27_109AddendStage1Output);

    MB_D_FF_Float_27_109_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF27_109AddendStage1Output, mb_D_FF27_109AddendStage2Output);

    MB_D_FF_Float_Multiplier10_Input1_82_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder27_Output_109, mb_D_FFMultiplier10_Input1_82_0Output);

    MB_D_FF_Float_82_110_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier10_Input1_82_0Output, mb_D_FF82_110MultiplicandStage1Output);

    MB_D_FF_Float_82_110_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF82_110MultiplicandStage1Output, mb_D_FF82_110MultiplicandStage2Output);

    Multiplier_Float_82: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF82_110MultiplicandStage2Output, mb_D_FF82_110MultiplierStage2Output, Multiplier82_Output_110);

    MB_D_FF_Float_Multiplier10_Input2_82_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier79_Output_106, mb_D_FFMultiplier10_Input2_82_0Output);

    MB_D_FF_Float_82_110_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier10_Input2_82_0Output, mb_D_FF82_110MultiplierStage1Output);

    MB_D_FF_Float_82_110_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF82_110MultiplierStage1Output, mb_D_FF82_110MultiplierStage2Output);

    MBRightSHR_Float_83_Input1111: entity work.MBRightSHR(rtl)
    GENERIC MAP (142, NumberOfBits)
    PORT MAP (clk, rst, Multiplier83Weight, mbRightSHR83_Input1_111Output);

    MB_D_FF_Float_83_111_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR83_Input1_111Output, Multiplier83WeightOutput);

    InputIEEE_Float_83_111: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier83WeightOutput, flopocoMultiplier83WeightOutput);

    MB_D_FF_Float_83_111_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier83WeightOutput, flopocoMultiplier83WeightInput);

    Multiplier_Float_83: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier83WeightInput, mb_D_FF83_111MultiplierStage2Output, Multiplier83_Output_111);

    MBRightSHR_Float_83_Input2_111: entity work.MBRightSHR(rtl)
    GENERIC MAP (142, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR83_Input2_111Input, mbRightSHR83_Input2_111Output);

    MB_D_FF_Float_83_111_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR83_Input2_111Output, mb_D_FF83_111MultiplierStage1Output);

    MB_D_FF_Float_83_111_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF83_111MultiplierStage1Output, mb_D_FF83_111MultiplierStage2Output);

    MBRightSHR_Float_84_Input1112: entity work.MBRightSHR(rtl)
    GENERIC MAP (142, NumberOfBits)
    PORT MAP (clk, rst, Multiplier84Weight, mbRightSHR84_Input1_112Output);

    MB_D_FF_Float_84_112_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR84_Input1_112Output, Multiplier84WeightOutput);

    InputIEEE_Float_84_112: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier84WeightOutput, flopocoMultiplier84WeightOutput);

    MB_D_FF_Float_84_112_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier84WeightOutput, flopocoMultiplier84WeightInput);

    Multiplier_Float_84: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier84WeightInput, mb_D_FF84_112MultiplierStage2Output, Multiplier84_Output_112);

    MBRightSHR_Float_84_Input2_112: entity work.MBRightSHR(rtl)
    GENERIC MAP (142, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR84_Input2_112Input, mbRightSHR84_Input2_112Output);

    MB_D_FF_Float_84_112_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR84_Input2_112Output, mb_D_FF84_112MultiplierStage1Output);

    MB_D_FF_Float_84_112_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF84_112MultiplierStage1Output, mb_D_FF84_112MultiplierStage2Output);

    MB_D_FF_Float_Adder10_Input1_28_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier84_Output_112, mb_D_FFAdder10_Input1_28_0Output);

    MB_D_FF_Float_28_113_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder10_Input1_28_0Output, mb_D_FF28_113AugendStage1Output);

    MB_D_FF_Float_28_113_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF28_113AugendStage1Output, mb_D_FF28_113AugendStage2Output);

    Adder_Float_28: entity work.FPAdd_7_24_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF28_113AugendStage2Output, mb_D_FF28_113AddendStage2Output, Adder28_Output_113);

    MB_D_FF_Float_Adder10_Input2_28_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier83_Output_111, mb_D_FFAdder10_Input2_28_0Output);

    MB_D_FF_Float_28_113_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder10_Input2_28_0Output, mb_D_FF28_113AddendStage1Output);

    MB_D_FF_Float_28_113_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF28_113AddendStage1Output, mb_D_FF28_113AddendStage2Output);

    MB_D_FF_Float_Multiplier9_Input1_85_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder28_Output_113, mb_D_FFMultiplier9_Input1_85_0Output);

    MB_D_FF_Float_85_114_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier9_Input1_85_0Output, mb_D_FF85_114MultiplicandStage1Output);

    MB_D_FF_Float_85_114_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF85_114MultiplicandStage1Output, mb_D_FF85_114MultiplicandStage2Output);

    Multiplier_Float_85: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF85_114MultiplicandStage2Output, mb_D_FF85_114MultiplierStage2Output, Multiplier85_Output_114);

    MB_D_FF_Float_Multiplier9_Input2_85_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier82_Output_110, mb_D_FFMultiplier9_Input2_85_0Output);

    MB_D_FF_Float_85_114_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier9_Input2_85_0Output, mb_D_FF85_114MultiplierStage1Output);

    MB_D_FF_Float_85_114_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF85_114MultiplierStage1Output, mb_D_FF85_114MultiplierStage2Output);

    MBRightSHR_Float_86_Input1115: entity work.MBRightSHR(rtl)
    GENERIC MAP (154, NumberOfBits)
    PORT MAP (clk, rst, Multiplier86Weight, mbRightSHR86_Input1_115Output);

    MB_D_FF_Float_86_115_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR86_Input1_115Output, Multiplier86WeightOutput);

    InputIEEE_Float_86_115: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier86WeightOutput, flopocoMultiplier86WeightOutput);

    MB_D_FF_Float_86_115_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier86WeightOutput, flopocoMultiplier86WeightInput);

    Multiplier_Float_86: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier86WeightInput, mb_D_FF86_115MultiplierStage2Output, Multiplier86_Output_115);

    MBRightSHR_Float_86_Input2_115: entity work.MBRightSHR(rtl)
    GENERIC MAP (154, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR86_Input2_115Input, mbRightSHR86_Input2_115Output);

    MB_D_FF_Float_86_115_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR86_Input2_115Output, mb_D_FF86_115MultiplierStage1Output);

    MB_D_FF_Float_86_115_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF86_115MultiplierStage1Output, mb_D_FF86_115MultiplierStage2Output);

    MBRightSHR_Float_87_Input1116: entity work.MBRightSHR(rtl)
    GENERIC MAP (154, NumberOfBits)
    PORT MAP (clk, rst, Multiplier87Weight, mbRightSHR87_Input1_116Output);

    MB_D_FF_Float_87_116_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR87_Input1_116Output, Multiplier87WeightOutput);

    InputIEEE_Float_87_116: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier87WeightOutput, flopocoMultiplier87WeightOutput);

    MB_D_FF_Float_87_116_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier87WeightOutput, flopocoMultiplier87WeightInput);

    Multiplier_Float_87: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier87WeightInput, mb_D_FF87_116MultiplierStage2Output, Multiplier87_Output_116);

    MBRightSHR_Float_87_Input2_116: entity work.MBRightSHR(rtl)
    GENERIC MAP (154, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR87_Input2_116Input, mbRightSHR87_Input2_116Output);

    MB_D_FF_Float_87_116_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR87_Input2_116Output, mb_D_FF87_116MultiplierStage1Output);

    MB_D_FF_Float_87_116_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF87_116MultiplierStage1Output, mb_D_FF87_116MultiplierStage2Output);

    MB_D_FF_Float_Adder9_Input1_29_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier87_Output_116, mb_D_FFAdder9_Input1_29_0Output);

    MB_D_FF_Float_29_117_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder9_Input1_29_0Output, mb_D_FF29_117AugendStage1Output);

    MB_D_FF_Float_29_117_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF29_117AugendStage1Output, mb_D_FF29_117AugendStage2Output);

    Adder_Float_29: entity work.FPAdd_7_24_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF29_117AugendStage2Output, mb_D_FF29_117AddendStage2Output, Adder29_Output_117);

    MB_D_FF_Float_Adder9_Input2_29_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier86_Output_115, mb_D_FFAdder9_Input2_29_0Output);

    MB_D_FF_Float_29_117_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder9_Input2_29_0Output, mb_D_FF29_117AddendStage1Output);

    MB_D_FF_Float_29_117_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF29_117AddendStage1Output, mb_D_FF29_117AddendStage2Output);

    MB_D_FF_Float_Multiplier8_Input1_88_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder29_Output_117, mb_D_FFMultiplier8_Input1_88_0Output);

    MB_D_FF_Float_88_118_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier8_Input1_88_0Output, mb_D_FF88_118MultiplicandStage1Output);

    MB_D_FF_Float_88_118_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF88_118MultiplicandStage1Output, mb_D_FF88_118MultiplicandStage2Output);

    Multiplier_Float_88: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF88_118MultiplicandStage2Output, mb_D_FF88_118MultiplierStage2Output, Multiplier88_Output_118);

    MB_D_FF_Float_Multiplier8_Input2_88_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier85_Output_114, mb_D_FFMultiplier8_Input2_88_0Output);

    MB_D_FF_Float_88_118_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier8_Input2_88_0Output, mb_D_FF88_118MultiplierStage1Output);

    MB_D_FF_Float_88_118_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF88_118MultiplierStage1Output, mb_D_FF88_118MultiplierStage2Output);

    MBRightSHR_Float_89_Input1119: entity work.MBRightSHR(rtl)
    GENERIC MAP (166, NumberOfBits)
    PORT MAP (clk, rst, Multiplier89Weight, mbRightSHR89_Input1_119Output);

    MB_D_FF_Float_89_119_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR89_Input1_119Output, Multiplier89WeightOutput);

    InputIEEE_Float_89_119: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier89WeightOutput, flopocoMultiplier89WeightOutput);

    MB_D_FF_Float_89_119_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier89WeightOutput, flopocoMultiplier89WeightInput);

    Multiplier_Float_89: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier89WeightInput, mb_D_FF89_119MultiplierStage2Output, Multiplier89_Output_119);

    MBRightSHR_Float_89_Input2_119: entity work.MBRightSHR(rtl)
    GENERIC MAP (166, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR89_Input2_119Input, mbRightSHR89_Input2_119Output);

    MB_D_FF_Float_89_119_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR89_Input2_119Output, mb_D_FF89_119MultiplierStage1Output);

    MB_D_FF_Float_89_119_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF89_119MultiplierStage1Output, mb_D_FF89_119MultiplierStage2Output);

    MBRightSHR_Float_90_Input1120: entity work.MBRightSHR(rtl)
    GENERIC MAP (166, NumberOfBits)
    PORT MAP (clk, rst, Multiplier90Weight, mbRightSHR90_Input1_120Output);

    MB_D_FF_Float_90_120_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR90_Input1_120Output, Multiplier90WeightOutput);

    InputIEEE_Float_90_120: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier90WeightOutput, flopocoMultiplier90WeightOutput);

    MB_D_FF_Float_90_120_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier90WeightOutput, flopocoMultiplier90WeightInput);

    Multiplier_Float_90: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier90WeightInput, mb_D_FF90_120MultiplierStage2Output, Multiplier90_Output_120);

    MBRightSHR_Float_90_Input2_120: entity work.MBRightSHR(rtl)
    GENERIC MAP (166, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR90_Input2_120Input, mbRightSHR90_Input2_120Output);

    MB_D_FF_Float_90_120_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR90_Input2_120Output, mb_D_FF90_120MultiplierStage1Output);

    MB_D_FF_Float_90_120_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF90_120MultiplierStage1Output, mb_D_FF90_120MultiplierStage2Output);

    MB_D_FF_Float_Adder8_Input1_30_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier90_Output_120, mb_D_FFAdder8_Input1_30_0Output);

    MB_D_FF_Float_30_121_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder8_Input1_30_0Output, mb_D_FF30_121AugendStage1Output);

    MB_D_FF_Float_30_121_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF30_121AugendStage1Output, mb_D_FF30_121AugendStage2Output);

    Adder_Float_30: entity work.FPAdd_7_24_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF30_121AugendStage2Output, mb_D_FF30_121AddendStage2Output, Adder30_Output_121);

    MB_D_FF_Float_Adder8_Input2_30_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier89_Output_119, mb_D_FFAdder8_Input2_30_0Output);

    MB_D_FF_Float_30_121_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder8_Input2_30_0Output, mb_D_FF30_121AddendStage1Output);

    MB_D_FF_Float_30_121_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF30_121AddendStage1Output, mb_D_FF30_121AddendStage2Output);

    MB_D_FF_Float_Multiplier7_Input1_91_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder30_Output_121, mb_D_FFMultiplier7_Input1_91_0Output);

    MB_D_FF_Float_91_122_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier7_Input1_91_0Output, mb_D_FF91_122MultiplicandStage1Output);

    MB_D_FF_Float_91_122_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF91_122MultiplicandStage1Output, mb_D_FF91_122MultiplicandStage2Output);

    Multiplier_Float_91: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF91_122MultiplicandStage2Output, mb_D_FF91_122MultiplierStage2Output, Multiplier91_Output_122);

    MB_D_FF_Float_Multiplier7_Input2_91_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier88_Output_118, mb_D_FFMultiplier7_Input2_91_0Output);

    MB_D_FF_Float_91_122_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier7_Input2_91_0Output, mb_D_FF91_122MultiplierStage1Output);

    MB_D_FF_Float_91_122_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF91_122MultiplierStage1Output, mb_D_FF91_122MultiplierStage2Output);

    MBRightSHR_Float_92_Input1123: entity work.MBRightSHR(rtl)
    GENERIC MAP (178, NumberOfBits)
    PORT MAP (clk, rst, Multiplier92Weight, mbRightSHR92_Input1_123Output);

    MB_D_FF_Float_92_123_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR92_Input1_123Output, Multiplier92WeightOutput);

    InputIEEE_Float_92_123: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier92WeightOutput, flopocoMultiplier92WeightOutput);

    MB_D_FF_Float_92_123_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier92WeightOutput, flopocoMultiplier92WeightInput);

    Multiplier_Float_92: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier92WeightInput, mb_D_FF92_123MultiplierStage2Output, Multiplier92_Output_123);

    MBRightSHR_Float_92_Input2_123: entity work.MBRightSHR(rtl)
    GENERIC MAP (178, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR92_Input2_123Input, mbRightSHR92_Input2_123Output);

    MB_D_FF_Float_92_123_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR92_Input2_123Output, mb_D_FF92_123MultiplierStage1Output);

    MB_D_FF_Float_92_123_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF92_123MultiplierStage1Output, mb_D_FF92_123MultiplierStage2Output);

    MBRightSHR_Float_93_Input1124: entity work.MBRightSHR(rtl)
    GENERIC MAP (178, NumberOfBits)
    PORT MAP (clk, rst, Multiplier93Weight, mbRightSHR93_Input1_124Output);

    MB_D_FF_Float_93_124_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR93_Input1_124Output, Multiplier93WeightOutput);

    InputIEEE_Float_93_124: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier93WeightOutput, flopocoMultiplier93WeightOutput);

    MB_D_FF_Float_93_124_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier93WeightOutput, flopocoMultiplier93WeightInput);

    Multiplier_Float_93: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier93WeightInput, mb_D_FF93_124MultiplierStage2Output, Multiplier93_Output_124);

    MBRightSHR_Float_93_Input2_124: entity work.MBRightSHR(rtl)
    GENERIC MAP (178, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR93_Input2_124Input, mbRightSHR93_Input2_124Output);

    MB_D_FF_Float_93_124_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR93_Input2_124Output, mb_D_FF93_124MultiplierStage1Output);

    MB_D_FF_Float_93_124_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF93_124MultiplierStage1Output, mb_D_FF93_124MultiplierStage2Output);

    MB_D_FF_Float_Adder7_Input1_31_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier93_Output_124, mb_D_FFAdder7_Input1_31_0Output);

    MB_D_FF_Float_31_125_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder7_Input1_31_0Output, mb_D_FF31_125AugendStage1Output);

    MB_D_FF_Float_31_125_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF31_125AugendStage1Output, mb_D_FF31_125AugendStage2Output);

    Adder_Float_31: entity work.FPAdd_7_24_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF31_125AugendStage2Output, mb_D_FF31_125AddendStage2Output, Adder31_Output_125);

    MB_D_FF_Float_Adder7_Input2_31_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier92_Output_123, mb_D_FFAdder7_Input2_31_0Output);

    MB_D_FF_Float_31_125_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder7_Input2_31_0Output, mb_D_FF31_125AddendStage1Output);

    MB_D_FF_Float_31_125_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF31_125AddendStage1Output, mb_D_FF31_125AddendStage2Output);

    MB_D_FF_Float_Multiplier6_Input1_94_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder31_Output_125, mb_D_FFMultiplier6_Input1_94_0Output);

    MB_D_FF_Float_94_126_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier6_Input1_94_0Output, mb_D_FF94_126MultiplicandStage1Output);

    MB_D_FF_Float_94_126_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF94_126MultiplicandStage1Output, mb_D_FF94_126MultiplicandStage2Output);

    Multiplier_Float_94: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF94_126MultiplicandStage2Output, mb_D_FF94_126MultiplierStage2Output, Multiplier94_Output_126);

    MB_D_FF_Float_Multiplier6_Input2_94_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier91_Output_122, mb_D_FFMultiplier6_Input2_94_0Output);

    MB_D_FF_Float_94_126_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier6_Input2_94_0Output, mb_D_FF94_126MultiplierStage1Output);

    MB_D_FF_Float_94_126_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF94_126MultiplierStage1Output, mb_D_FF94_126MultiplierStage2Output);

    MBRightSHR_Float_95_Input1127: entity work.MBRightSHR(rtl)
    GENERIC MAP (190, NumberOfBits)
    PORT MAP (clk, rst, Multiplier95Weight, mbRightSHR95_Input1_127Output);

    MB_D_FF_Float_95_127_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR95_Input1_127Output, Multiplier95WeightOutput);

    InputIEEE_Float_95_127: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier95WeightOutput, flopocoMultiplier95WeightOutput);

    MB_D_FF_Float_95_127_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier95WeightOutput, flopocoMultiplier95WeightInput);

    Multiplier_Float_95: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier95WeightInput, mb_D_FF95_127MultiplierStage2Output, Multiplier95_Output_127);

    MBRightSHR_Float_95_Input2_127: entity work.MBRightSHR(rtl)
    GENERIC MAP (190, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR95_Input2_127Input, mbRightSHR95_Input2_127Output);

    MB_D_FF_Float_95_127_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR95_Input2_127Output, mb_D_FF95_127MultiplierStage1Output);

    MB_D_FF_Float_95_127_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF95_127MultiplierStage1Output, mb_D_FF95_127MultiplierStage2Output);

    MBRightSHR_Float_96_Input1128: entity work.MBRightSHR(rtl)
    GENERIC MAP (190, NumberOfBits)
    PORT MAP (clk, rst, Multiplier96Weight, mbRightSHR96_Input1_128Output);

    MB_D_FF_Float_96_128_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR96_Input1_128Output, Multiplier96WeightOutput);

    InputIEEE_Float_96_128: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier96WeightOutput, flopocoMultiplier96WeightOutput);

    MB_D_FF_Float_96_128_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier96WeightOutput, flopocoMultiplier96WeightInput);

    Multiplier_Float_96: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier96WeightInput, mb_D_FF96_128MultiplierStage2Output, Multiplier96_Output_128);

    MBRightSHR_Float_96_Input2_128: entity work.MBRightSHR(rtl)
    GENERIC MAP (190, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR96_Input2_128Input, mbRightSHR96_Input2_128Output);

    MB_D_FF_Float_96_128_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR96_Input2_128Output, mb_D_FF96_128MultiplierStage1Output);

    MB_D_FF_Float_96_128_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF96_128MultiplierStage1Output, mb_D_FF96_128MultiplierStage2Output);

    MB_D_FF_Float_Adder6_Input1_32_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier96_Output_128, mb_D_FFAdder6_Input1_32_0Output);

    MB_D_FF_Float_32_129_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder6_Input1_32_0Output, mb_D_FF32_129AugendStage1Output);

    MB_D_FF_Float_32_129_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF32_129AugendStage1Output, mb_D_FF32_129AugendStage2Output);

    Adder_Float_32: entity work.FPAdd_7_24_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF32_129AugendStage2Output, mb_D_FF32_129AddendStage2Output, Adder32_Output_129);

    MB_D_FF_Float_Adder6_Input2_32_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier95_Output_127, mb_D_FFAdder6_Input2_32_0Output);

    MB_D_FF_Float_32_129_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder6_Input2_32_0Output, mb_D_FF32_129AddendStage1Output);

    MB_D_FF_Float_32_129_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF32_129AddendStage1Output, mb_D_FF32_129AddendStage2Output);

    MB_D_FF_Float_Multiplier5_Input1_97_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder32_Output_129, mb_D_FFMultiplier5_Input1_97_0Output);

    MB_D_FF_Float_97_130_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier5_Input1_97_0Output, mb_D_FF97_130MultiplicandStage1Output);

    MB_D_FF_Float_97_130_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF97_130MultiplicandStage1Output, mb_D_FF97_130MultiplicandStage2Output);

    Multiplier_Float_97: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF97_130MultiplicandStage2Output, mb_D_FF97_130MultiplierStage2Output, Multiplier97_Output_130);

    MB_D_FF_Float_Multiplier5_Input2_97_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier94_Output_126, mb_D_FFMultiplier5_Input2_97_0Output);

    MB_D_FF_Float_97_130_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier5_Input2_97_0Output, mb_D_FF97_130MultiplierStage1Output);

    MB_D_FF_Float_97_130_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF97_130MultiplierStage1Output, mb_D_FF97_130MultiplierStage2Output);

    MBRightSHR_Float_98_Input1131: entity work.MBRightSHR(rtl)
    GENERIC MAP (202, NumberOfBits)
    PORT MAP (clk, rst, Multiplier98Weight, mbRightSHR98_Input1_131Output);

    MB_D_FF_Float_98_131_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR98_Input1_131Output, Multiplier98WeightOutput);

    InputIEEE_Float_98_131: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier98WeightOutput, flopocoMultiplier98WeightOutput);

    MB_D_FF_Float_98_131_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier98WeightOutput, flopocoMultiplier98WeightInput);

    Multiplier_Float_98: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier98WeightInput, mb_D_FF98_131MultiplierStage2Output, Multiplier98_Output_131);

    MBRightSHR_Float_98_Input2_131: entity work.MBRightSHR(rtl)
    GENERIC MAP (202, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR98_Input2_131Input, mbRightSHR98_Input2_131Output);

    MB_D_FF_Float_98_131_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR98_Input2_131Output, mb_D_FF98_131MultiplierStage1Output);

    MB_D_FF_Float_98_131_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF98_131MultiplierStage1Output, mb_D_FF98_131MultiplierStage2Output);

    MBRightSHR_Float_99_Input1132: entity work.MBRightSHR(rtl)
    GENERIC MAP (202, NumberOfBits)
    PORT MAP (clk, rst, Multiplier99Weight, mbRightSHR99_Input1_132Output);

    MB_D_FF_Float_99_132_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR99_Input1_132Output, Multiplier99WeightOutput);

    InputIEEE_Float_99_132: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier99WeightOutput, flopocoMultiplier99WeightOutput);

    MB_D_FF_Float_99_132_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier99WeightOutput, flopocoMultiplier99WeightInput);

    Multiplier_Float_99: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, flopocoMultiplier99WeightInput, mb_D_FF99_132MultiplierStage2Output, Multiplier99_Output_132);

    MBRightSHR_Float_99_Input2_132: entity work.MBRightSHR(rtl)
    GENERIC MAP (202, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR99_Input2_132Input, mbRightSHR99_Input2_132Output);

    MB_D_FF_Float_99_132_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR99_Input2_132Output, mb_D_FF99_132MultiplierStage1Output);

    MB_D_FF_Float_99_132_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF99_132MultiplierStage1Output, mb_D_FF99_132MultiplierStage2Output);

    MB_D_FF_Float_Adder5_Input1_33_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier99_Output_132, mb_D_FFAdder5_Input1_33_0Output);

    MB_D_FF_Float_33_133_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder5_Input1_33_0Output, mb_D_FF33_133AugendStage1Output);

    MB_D_FF_Float_33_133_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF33_133AugendStage1Output, mb_D_FF33_133AugendStage2Output);

    Adder_Float_33: entity work.FPAdd_7_24_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF33_133AugendStage2Output, mb_D_FF33_133AddendStage2Output, Adder33_Output_133);

    MB_D_FF_Float_Adder5_Input2_33_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier98_Output_131, mb_D_FFAdder5_Input2_33_0Output);

    MB_D_FF_Float_33_133_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder5_Input2_33_0Output, mb_D_FF33_133AddendStage1Output);

    MB_D_FF_Float_33_133_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF33_133AddendStage1Output, mb_D_FF33_133AddendStage2Output);

    MB_D_FF_Float_Multiplier4_Input1_100_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder33_Output_133, mb_D_FFMultiplier4_Input1_100_0Output);

    MB_D_FF_Float_100_134_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier4_Input1_100_0Output, mb_D_FF100_134MultiplicandStage1Output);

    MB_D_FF_Float_100_134_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF100_134MultiplicandStage1Output, mb_D_FF100_134MultiplicandStage2Output);

    Multiplier_Float_100: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF100_134MultiplicandStage2Output, mb_D_FF100_134MultiplierStage2Output, Multiplier100_Output_134);

    MB_D_FF_Float_Multiplier4_Input2_100_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier97_Output_130, mb_D_FFMultiplier4_Input2_100_0Output);

    MB_D_FF_Float_100_134_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier4_Input2_100_0Output, mb_D_FF100_134MultiplierStage1Output);

    MB_D_FF_Float_100_134_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF100_134MultiplierStage1Output, mb_D_FF100_134MultiplierStage2Output);

    MB_D_FF_Float_Multiplier3_101_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier100_Output_134, mb_D_FFMultiplier3_101_0Output);

    MB_D_FF_Float_101_135_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier3_101_0Output, mb_D_FF101_135MultiplierStage1Output);

    MB_D_FF_Float_101_135_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF101_135MultiplierStage1Output, mb_D_FF101_135MultiplierStage2Output);

    Multiplier_Float_101: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF101_135MultiplierStage2Output, mb_D_FF101_135MultiplicandStage2Output, Multiplier101_Output_135);

    MBRightSHR_Float_101_135: entity work.MBRightSHR(rtl)
    GENERIC MAP (238, NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR101_135Input, mbRightSHR101_135Output);

    MB_D_FF_Float_101_135_MultiplicandStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mbRightSHR101_135Output, mb_D_FF101_135MultiplicandStage1Output);

    MB_D_FF_Float_101_135_MultiplicandStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF101_135MultiplicandStage1Output, mb_D_FF101_135MultiplicandStage2Output);

    MB_D_FF_Float_Multiplier2_102_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier101_Output_135, mb_D_FFMultiplier2_102_0Output);

    MB_D_FF_Float_102_136_MultiplierStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFMultiplier2_102_0Output, mb_D_FF102_136MultiplierStage1Output);

    MB_D_FF_Float_102_136_MultiplierStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF102_136MultiplierStage1Output, mb_D_FF102_136MultiplierStage2Output);

    Multiplier_Float_102: entity work.FPMult_7_24_7_24_7_24_uid2_Freq800_uid3(arch)
    PORT MAP (clk, mb_D_FF102_136MultiplierStage2Output, flopocoMultiplier102WeightInput, Multiplier102_Output_136);

    MBRightSHR_Float_102_136: entity work.MBRightSHR(rtl)
    GENERIC MAP (250, NumberOfBits)
    PORT MAP (clk, rst, Multiplier102Weight, mbRightSHR102_136Output);

    MB_D_FF_Float_102_136_ConverterInput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits)
    PORT MAP (clk, rst, mbRightSHR102_136Output, Multiplier102WeightOutput);

    InputIEEE_Float_102_136: entity work.InputIEEE_7_24_to_7_24(arch)
        PORT MAP (clk, Multiplier102WeightOutput, flopocoMultiplier102WeightOutput);

    MB_D_FF_Float_102_136_ConverterOutput: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, flopocoMultiplier102WeightOutput, flopocoMultiplier102WeightInput);

    MB_D_FF_Float_Adder1_Input1_34_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier102_Output_136, mb_D_FFAdder1_Input1_34_0Output);

    MB_D_FF_Float_34_137_AugendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder1_Input1_34_0Output, mb_D_FF34_137AugendStage1Output);

    MB_D_FF_Float_34_137_AugendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF34_137AugendStage1Output, mb_D_FF34_137AugendStage2Output);

    Adder_Float_34: entity work.FPAdd_7_24_Freq800_uid2(arch)
    PORT MAP (clk, mb_D_FF34_137AugendStage2Output, mb_D_FF34_137AddendStage2Output, Adder34_Output_137);

    MB_D_FF_Float_Adder1_Input2_34_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Multiplier53_Output_71, mb_D_FFAdder1_Input2_34_0Output);

    MB_D_FF_Float_34_137_AddendStage1Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FFAdder1_Input2_34_0Output, mb_D_FF34_137AddendStage1Output);

    MB_D_FF_Float_34_137_AddendStage2Register: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, mb_D_FF34_137AddendStage1Output, mb_D_FF34_137AddendStage2Output);

    MB_D_FF_Float_Adder1_Output_34_0: entity work.MB_D_FF(rtl)
    GENERIC MAP (NumberOfBits+FlopocoBits)
    PORT MAP (clk, rst, Adder34_Output_137, mb_D_FFAdder1_Output_34_0Output);

    vout <= mb_D_FFAdder1_Output_34_0Output;
 
END ARCHITECTURE;

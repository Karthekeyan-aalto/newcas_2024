library ieee; 
library ieee_proposed; 
use ieee.std_logic_1164.all; 
use ieee.numeric_std.all; 
use std.textio.all; 
use ieee_proposed.fixed_pkg.all; 
use ieee_proposed.fixed_float_types.all; 
USE ieee_proposed.float_pkg.all; 
 
entity PCSystem is 
 
generic(mantissaBits : integer := 15; exponentBits : integer := 5);
port( 
v1 : in float (5 DOWNTO -14);
v2 : in float (5 DOWNTO -14);
v3 : in float (5 DOWNTO -14);
v4 : in float (5 DOWNTO -14);
v5 : in float (5 DOWNTO -14);
v6 : in float (5 DOWNTO -14);
v7 : in float (5 DOWNTO -14);
v8 : in float (5 DOWNTO -14);
v9 : in float (5 DOWNTO -14);
v10 : in float (5 DOWNTO -14);
v11 : in float (5 DOWNTO -14);
v12 : in float (5 DOWNTO -14);
v13 : in float (5 DOWNTO -14);
v14 : in float (5 DOWNTO -14);
v15 : in float (5 DOWNTO -14);
v16 : in float (5 DOWNTO -14);
vb1 : in float (5 DOWNTO -14);
vb2 : in float (5 DOWNTO -14);
vb3 : in float (5 DOWNTO -14);
vb4 : in float (5 DOWNTO -14);
vb5 : in float (5 DOWNTO -14);
vb6 : in float (5 DOWNTO -14);
vb7 : in float (5 DOWNTO -14);
vb8 : in float (5 DOWNTO -14);
vb9 : in float (5 DOWNTO -14);
vb10 : in float (5 DOWNTO -14);
vb11 : in float (5 DOWNTO -14);
vb12 : in float (5 DOWNTO -14);
vb13 : in float (5 DOWNTO -14);
vb14 : in float (5 DOWNTO -14);
vb15 : in float (5 DOWNTO -14);
vb16 : in float (5 DOWNTO -14);
vout : out float (5 DOWNTO -14)); 
 
end PCSystem; 

architecture rtl of PCSystem is 
 
Signal ProductNode_Float0weight : float ( 5 downto -14 ) := to_float (0.848299,5,14);

Signal ProductNode_Float0Output_0: float (5 downto -14);
Signal ProductNode_Float1weight : float ( 5 downto -14 ) := to_float (0.895308,5,14);

Signal ProductNode_Float1Output_1: float (5 downto -14);
Signal ProductNode_Float2weight : float ( 5 downto -14 ) := to_float (0.842608,5,14);

Signal ProductNode_Float2Output_2: float (5 downto -14);
Signal SumNode_Float0Output_3: float (5 downto -14);
Signal ProductNode_Float3Output_4: float (5 downto -14);
Signal ProductNode_Float4weight : float ( 5 downto -14 ) := to_float (0.870697,5,14);

Signal ProductNode_Float4Output_5: float (5 downto -14);
Signal ProductNode_Float5weight : float ( 5 downto -14 ) := to_float (0.945793,5,14);

Signal ProductNode_Float5Output_6: float (5 downto -14);
Signal ProductNode_Float6weight : float ( 5 downto -14 ) := to_float (0.954870,5,14);

Signal ProductNode_Float6Output_7: float (5 downto -14);
Signal ProductNode_Float7weight : float ( 5 downto -14 ) := to_float (0.870404,5,14);

Signal ProductNode_Float7Output_8: float (5 downto -14);
Signal ProductNode_Float8weight : float ( 5 downto -14 ) := to_float (0.780732,5,14);

Signal ProductNode_Float8Output_9: float (5 downto -14);
Signal ProductNode_Float9weight : float ( 5 downto -14 ) := to_float (0.810846,5,14);

Signal ProductNode_Float9Output_10: float (5 downto -14);
Signal SumNode_Float1Output_11: float (5 downto -14);
Signal ProductNode_Float10Output_12: float (5 downto -14);
Signal ProductNode_Float11weight : float ( 5 downto -14 ) := to_float (0.991361,5,14);

Signal ProductNode_Float11Output_13: float (5 downto -14);
Signal ProductNode_Float12weight : float ( 5 downto -14 ) := to_float (0.669241,5,14);

Signal ProductNode_Float12Output_14: float (5 downto -14);
Signal ProductNode_Float13weight : float ( 5 downto -14 ) := to_float (0.971580,5,14);

Signal ProductNode_Float13Output_15: float (5 downto -14);
Signal SumNode_Float2Output_16: float (5 downto -14);
Signal ProductNode_Float14Output_17: float (5 downto -14);
Signal ProductNode_Float15weight : float ( 5 downto -14 ) := to_float (0.870697,5,14);

Signal ProductNode_Float15Output_18: float (5 downto -14);
Signal ProductNode_Float16weight : float ( 5 downto -14 ) := to_float (0.753690,5,14);

Signal ProductNode_Float16Output_19: float (5 downto -14);
Signal ProductNode_Float17weight : float ( 5 downto -14 ) := to_float (0.774480,5,14);

Signal ProductNode_Float17Output_20: float (5 downto -14);
Signal ProductNode_Float18weight : float ( 5 downto -14 ) := to_float (0.870404,5,14);

Signal ProductNode_Float18Output_21: float (5 downto -14);
Signal ProductNode_Float19weight : float ( 5 downto -14 ) := to_float (0.933776,5,14);

Signal ProductNode_Float19Output_22: float (5 downto -14);
Signal ProductNode_Float20weight : float ( 5 downto -14 ) := to_float (0.660973,5,14);

Signal ProductNode_Float20Output_23: float (5 downto -14);
Signal SumNode_Float3Output_24: float (5 downto -14);
Signal ProductNode_Float21Output_25: float (5 downto -14);
Signal ProductNode_Float22weight : float ( 5 downto -14 ) := to_float (0.870239,5,14);

Signal ProductNode_Float22Output_26: float (5 downto -14);
Signal SumNode_Float4Output_27: float (5 downto -14);
Signal ProductNode_Float23Output_28: float (5 downto -14);
Signal ProductNode_Float24weight : float ( 5 downto -14 ) := to_float (0.944720,5,14);

Signal ProductNode_Float24Output_29: float (5 downto -14);
Signal ProductNode_Float25weight : float ( 5 downto -14 ) := to_float (0.890735,5,14);

Signal ProductNode_Float25Output_30: float (5 downto -14);
Signal ProductNode_Float26weight : float ( 5 downto -14 ) := to_float (0.689002,5,14);

Signal ProductNode_Float26Output_31: float (5 downto -14);
Signal ProductNode_Float27weight : float ( 5 downto -14 ) := to_float (0.966814,5,14);

Signal ProductNode_Float27Output_32: float (5 downto -14);
Signal SumNode_Float5Output_33: float (5 downto -14);
Signal ProductNode_Float28Output_34: float (5 downto -14);
Signal ProductNode_Float29weight : float ( 5 downto -14 ) := to_float (0.551341,5,14);

Signal ProductNode_Float29Output_35: float (5 downto -14);
Signal ProductNode_Float30weight : float ( 5 downto -14 ) := to_float (0.795357,5,14);

Signal ProductNode_Float30Output_36: float (5 downto -14);
Signal ProductNode_Float31weight : float ( 5 downto -14 ) := to_float (0.746308,5,14);

Signal ProductNode_Float31Output_37: float (5 downto -14);
Signal ProductNode_Float32weight : float ( 5 downto -14 ) := to_float (0.989597,5,14);

Signal ProductNode_Float32Output_38: float (5 downto -14);
Signal ProductNode_Float33weight : float ( 5 downto -14 ) := to_float (0.577708,5,14);

Signal ProductNode_Float33Output_39: float (5 downto -14);
Signal ProductNode_Float34weight : float ( 5 downto -14 ) := to_float (0.618274,5,14);

Signal ProductNode_Float34Output_40: float (5 downto -14);
Signal SumNode_Float6Output_41: float (5 downto -14);
Signal ProductNode_Float35Output_42: float (5 downto -14);
Signal ProductNode_Float36weight : float ( 5 downto -14 ) := to_float (0.952809,5,14);

Signal ProductNode_Float36Output_43: float (5 downto -14);
Signal ProductNode_Float37weight : float ( 5 downto -14 ) := to_float (0.495915,5,14);

Signal ProductNode_Float37Output_44: float (5 downto -14);
Signal ProductNode_Float38weight : float ( 5 downto -14 ) := to_float (0.993928,5,14);

Signal ProductNode_Float38Output_45: float (5 downto -14);
Signal SumNode_Float7Output_46: float (5 downto -14);
Signal ProductNode_Float39Output_47: float (5 downto -14);
Signal ProductNode_Float40weight : float ( 5 downto -14 ) := to_float (0.551341,5,14);

Signal ProductNode_Float40Output_48: float (5 downto -14);
Signal ProductNode_Float41weight : float ( 5 downto -14 ) := to_float (0.926235,5,14);

Signal ProductNode_Float41Output_49: float (5 downto -14);
Signal ProductNode_Float42weight : float ( 5 downto -14 ) := to_float (0.616494,5,14);

Signal ProductNode_Float42Output_50: float (5 downto -14);
Signal ProductNode_Float43weight : float ( 5 downto -14 ) := to_float (0.989597,5,14);

Signal ProductNode_Float43Output_51: float (5 downto -14);
Signal ProductNode_Float44weight : float ( 5 downto -14 ) := to_float (0.986786,5,14);

Signal ProductNode_Float44Output_52: float (5 downto -14);
Signal ProductNode_Float45weight : float ( 5 downto -14 ) := to_float (0.464416,5,14);

Signal ProductNode_Float45Output_53: float (5 downto -14);
Signal SumNode_Float8Output_54: float (5 downto -14);
Signal ProductNode_Float46Output_55: float (5 downto -14);
Signal ProductNode_Float47weight : float ( 5 downto -14 ) := to_float (0.770987,5,14);

Signal ProductNode_Float47Output_56: float (5 downto -14);
Signal SumNode_Float9Output_57: float (5 downto -14);
Signal ProductNode_Float48Output_58: float (5 downto -14);
Signal ProductNode_Float49weight : float ( 5 downto -14 ) := to_float (0.827729,5,14);

Signal ProductNode_Float49Output_59: float (5 downto -14);
Signal SumNode_Float10Output_60: float (5 downto -14);
Signal ProductNode_Float50Output_61: float (5 downto -14);
Signal ProductNode_Float51weight : float ( 5 downto -14 ) := to_float (0.986612,5,14);

Signal ProductNode_Float51Output_62: float (5 downto -14);
Signal ProductNode_Float52weight : float ( 5 downto -14 ) := to_float (0.848299,5,14);

Signal ProductNode_Float52Output_63: float (5 downto -14);
Signal ProductNode_Float53weight : float ( 5 downto -14 ) := to_float (0.562709,5,14);

Signal ProductNode_Float53Output_64: float (5 downto -14);
Signal ProductNode_Float54weight : float ( 5 downto -14 ) := to_float (0.988453,5,14);

Signal ProductNode_Float54Output_65: float (5 downto -14);
Signal SumNode_Float11Output_66: float (5 downto -14);
Signal ProductNode_Float55Output_67: float (5 downto -14);
Signal ProductNode_Float56weight : float ( 5 downto -14 ) := to_float (0.870697,5,14);

Signal ProductNode_Float56Output_68: float (5 downto -14);
Signal ProductNode_Float57weight : float ( 5 downto -14 ) := to_float (0.945793,5,14);

Signal ProductNode_Float57Output_69: float (5 downto -14);
Signal ProductNode_Float58weight : float ( 5 downto -14 ) := to_float (0.729204,5,14);

Signal ProductNode_Float58Output_70: float (5 downto -14);
Signal ProductNode_Float59weight : float ( 5 downto -14 ) := to_float (0.870404,5,14);

Signal ProductNode_Float59Output_71: float (5 downto -14);
Signal ProductNode_Float60weight : float ( 5 downto -14 ) := to_float (0.780732,5,14);

Signal ProductNode_Float60Output_72: float (5 downto -14);
Signal ProductNode_Float61weight : float ( 5 downto -14 ) := to_float (0.917308,5,14);

Signal ProductNode_Float61Output_73: float (5 downto -14);
Signal SumNode_Float12Output_74: float (5 downto -14);
Signal ProductNode_Float62Output_75: float (5 downto -14);
Signal ProductNode_Float63weight : float ( 5 downto -14 ) := to_float (0.979033,5,14);

Signal ProductNode_Float63Output_76: float (5 downto -14);
Signal ProductNode_Float64weight : float ( 5 downto -14 ) := to_float (0.453222,5,14);

Signal ProductNode_Float64Output_77: float (5 downto -14);
Signal ProductNode_Float65weight : float ( 5 downto -14 ) := to_float (0.996146,5,14);

Signal ProductNode_Float65Output_78: float (5 downto -14);
Signal SumNode_Float13Output_79: float (5 downto -14);
Signal ProductNode_Float66Output_80: float (5 downto -14);
Signal ProductNode_Float67weight : float ( 5 downto -14 ) := to_float (0.870697,5,14);

Signal ProductNode_Float67Output_81: float (5 downto -14);
Signal ProductNode_Float68weight : float ( 5 downto -14 ) := to_float (0.753690,5,14);

Signal ProductNode_Float68Output_82: float (5 downto -14);
Signal ProductNode_Float69weight : float ( 5 downto -14 ) := to_float (0.936763,5,14);

Signal ProductNode_Float69Output_83: float (5 downto -14);
Signal ProductNode_Float70weight : float ( 5 downto -14 ) := to_float (0.870404,5,14);

Signal ProductNode_Float70Output_84: float (5 downto -14);
Signal ProductNode_Float71weight : float ( 5 downto -14 ) := to_float (0.933776,5,14);

Signal ProductNode_Float71Output_85: float (5 downto -14);
Signal ProductNode_Float72weight : float ( 5 downto -14 ) := to_float (0.973389,5,14);

Signal ProductNode_Float72Output_86: float (5 downto -14);
Signal SumNode_Float14Output_87: float (5 downto -14);
Signal ProductNode_Float73Output_88: float (5 downto -14);
Signal ProductNode_Float74weight : float ( 5 downto -14 ) := to_float (0.818419,5,14);

Signal ProductNode_Float74Output_89: float (5 downto -14);
Signal SumNode_Float15Output_90: float (5 downto -14);
Signal ProductNode_Float75Output_91: float (5 downto -14);
Signal ProductNode_Float76weight : float ( 5 downto -14 ) := to_float (0.766253,5,14);

Signal ProductNode_Float76Output_92: float (5 downto -14);
Signal ProductNode_Float77weight : float ( 5 downto -14 ) := to_float (0.890735,5,14);

Signal ProductNode_Float77Output_93: float (5 downto -14);
Signal ProductNode_Float78weight : float ( 5 downto -14 ) := to_float (0.382644,5,14);

Signal ProductNode_Float78Output_94: float (5 downto -14);
Signal ProductNode_Float79weight : float ( 5 downto -14 ) := to_float (0.998354,5,14);

Signal ProductNode_Float79Output_95: float (5 downto -14);
Signal SumNode_Float16Output_96: float (5 downto -14);
Signal ProductNode_Float80Output_97: float (5 downto -14);
Signal ProductNode_Float81weight : float ( 5 downto -14 ) := to_float (0.551341,5,14);

Signal ProductNode_Float81Output_98: float (5 downto -14);
Signal ProductNode_Float82weight : float ( 5 downto -14 ) := to_float (0.795357,5,14);

Signal ProductNode_Float82Output_99: float (5 downto -14);
Signal ProductNode_Float83weight : float ( 5 downto -14 ) := to_float (0.948695,5,14);

Signal ProductNode_Float83Output_100: float (5 downto -14);
Signal ProductNode_Float84weight : float ( 5 downto -14 ) := to_float (0.989597,5,14);

Signal ProductNode_Float84Output_101: float (5 downto -14);
Signal ProductNode_Float85weight : float ( 5 downto -14 ) := to_float (0.577708,5,14);

Signal ProductNode_Float85Output_102: float (5 downto -14);
Signal ProductNode_Float86weight : float ( 5 downto -14 ) := to_float (0.981240,5,14);

Signal ProductNode_Float86Output_103: float (5 downto -14);
Signal SumNode_Float17Output_104: float (5 downto -14);
Signal ProductNode_Float87Output_105: float (5 downto -14);
Signal ProductNode_Float88weight : float ( 5 downto -14 ) := to_float (0.960334,5,14);

Signal ProductNode_Float88Output_106: float (5 downto -14);
Signal ProductNode_Float89weight : float ( 5 downto -14 ) := to_float (0.336149,5,14);

Signal ProductNode_Float89Output_107: float (5 downto -14);
Signal ProductNode_Float90weight : float ( 5 downto -14 ) := to_float (0.999140,5,14);

Signal ProductNode_Float90Output_108: float (5 downto -14);
Signal SumNode_Float18Output_109: float (5 downto -14);
Signal ProductNode_Float91Output_110: float (5 downto -14);
Signal ProductNode_Float92weight : float ( 5 downto -14 ) := to_float (0.551341,5,14);

Signal ProductNode_Float92Output_111: float (5 downto -14);
Signal ProductNode_Float93weight : float ( 5 downto -14 ) := to_float (0.926235,5,14);

Signal ProductNode_Float93Output_112: float (5 downto -14);
Signal ProductNode_Float94weight : float ( 5 downto -14 ) := to_float (0.981519,5,14);

Signal ProductNode_Float94Output_113: float (5 downto -14);
Signal ProductNode_Float95weight : float ( 5 downto -14 ) := to_float (0.989597,5,14);

Signal ProductNode_Float95Output_114: float (5 downto -14);
Signal ProductNode_Float96weight : float ( 5 downto -14 ) := to_float (0.986786,5,14);

Signal ProductNode_Float96Output_115: float (5 downto -14);
Signal ProductNode_Float97weight : float ( 5 downto -14 ) := to_float (0.995641,5,14);

Signal ProductNode_Float97Output_116: float (5 downto -14);
Signal SumNode_Float19Output_117: float (5 downto -14);
Signal ProductNode_Float98Output_118: float (5 downto -14);
Signal ProductNode_Float99weight : float ( 5 downto -14 ) := to_float (0.664315,5,14);

Signal ProductNode_Float99Output_119: float (5 downto -14);
Signal SumNode_Float20Output_120: float (5 downto -14);
Signal ProductNode_Float100Output_121: float (5 downto -14);
Signal ProductNode_Float101weight : float ( 5 downto -14 ) := to_float (0.634118,5,14);

Signal ProductNode_Float101Output_122: float (5 downto -14);
Signal SumNode_Float21Output_123: float (5 downto -14);
Signal ProductNode_Float102Output_124: float (5 downto -14);
Signal ProductNode_Float103weight : float ( 5 downto -14 ) := to_float (0.943120,5,14);

Signal ProductNode_Float103Output_125: float (5 downto -14);
Signal SumNode_Float22Output_126: float (5 downto -14);
Signal ProductNode_Float104Output_127: float (5 downto -14);
Signal ProductNode_Float105weight : float ( 5 downto -14 ) := to_float (0.970921,5,14);

Signal ProductNode_Float105Output_128: float (5 downto -14);
Signal ProductNode_Float106weight : float ( 5 downto -14 ) := to_float (0.672140,5,14);

Signal ProductNode_Float106Output_129: float (5 downto -14);
Signal SumNode_Float23Output_130: float (5 downto -14);
Signal ProductNode_Float107Output_131: float (5 downto -14);
Signal ProductNode_Float108weight : float ( 5 downto -14 ) := to_float (0.989270,5,14);

Signal ProductNode_Float108Output_132: float (5 downto -14);
Signal ProductNode_Float109weight : float ( 5 downto -14 ) := to_float (0.997554,5,14);

Signal ProductNode_Float109Output_133: float (5 downto -14);
Signal ProductNode_Float110weight : float ( 5 downto -14 ) := to_float (0.414069,5,14);

Signal ProductNode_Float110Output_134: float (5 downto -14);
Signal SumNode_Float24Output_135: float (5 downto -14);
Signal ProductNode_Float111Output_136: float (5 downto -14);
Signal ProductNode_Float112weight : float ( 5 downto -14 ) := to_float (0.853307,5,14);

Signal ProductNode_Float112Output_137: float (5 downto -14);
Signal ProductNode_Float113weight : float ( 5 downto -14 ) := to_float (0.886527,5,14);

Signal ProductNode_Float113Output_138: float (5 downto -14);
Signal SumNode_Float25Output_139: float (5 downto -14);
Signal ProductNode_Float114Output_140: float (5 downto -14);
Signal ProductNode_Float115weight : float ( 5 downto -14 ) := to_float (0.554692,5,14);

Signal ProductNode_Float115Output_141: float (5 downto -14);
Signal ProductNode_Float116weight : float ( 5 downto -14 ) := to_float (0.989739,5,14);

Signal ProductNode_Float116Output_142: float (5 downto -14);
Signal ProductNode_Float117weight : float ( 5 downto -14 ) := to_float (0.549861,5,14);

Signal ProductNode_Float117Output_143: float (5 downto -14);
Signal SumNode_Float26Output_144: float (5 downto -14);
Signal ProductNode_Float118Output_145: float (5 downto -14);
Signal SumNode_Float27Output_146: float (5 downto -14);
Signal ProductNode_Float119Output_147: float (5 downto -14);
Signal ProductNode_Float120weight : float ( 5 downto -14 ) := to_float (0.994862,5,14);

Signal ProductNode_Float120Output_148: float (5 downto -14);
Signal ProductNode_Float121weight : float ( 5 downto -14 ) := to_float (0.817897,5,14);

Signal ProductNode_Float121Output_149: float (5 downto -14);
Signal ProductNode_Float122weight : float ( 5 downto -14 ) := to_float (0.912886,5,14);

Signal ProductNode_Float122Output_150: float (5 downto -14);
Signal SumNode_Float28Output_151: float (5 downto -14);
Signal ProductNode_Float123Output_152: float (5 downto -14);
Signal ProductNode_Float124weight : float ( 5 downto -14 ) := to_float (0.976301,5,14);

Signal ProductNode_Float124Output_153: float (5 downto -14);
Signal ProductNode_Float125weight : float ( 5 downto -14 ) := to_float (0.988880,5,14);

Signal ProductNode_Float125Output_154: float (5 downto -14);
Signal ProductNode_Float126weight : float ( 5 downto -14 ) := to_float (0.558577,5,14);

Signal ProductNode_Float126Output_155: float (5 downto -14);
Signal SumNode_Float29Output_156: float (5 downto -14);
Signal ProductNode_Float127Output_157: float (5 downto -14);
Signal ProductNode_Float128weight : float ( 5 downto -14 ) := to_float (0.731617,5,14);

Signal ProductNode_Float128Output_158: float (5 downto -14);
Signal ProductNode_Float129weight : float ( 5 downto -14 ) := to_float (0.954043,5,14);

Signal ProductNode_Float129Output_159: float (5 downto -14);
Signal SumNode_Float30Output_160: float (5 downto -14);
Signal ProductNode_Float130Output_161: float (5 downto -14);
Signal ProductNode_Float131weight : float ( 5 downto -14 ) := to_float (0.646579,5,14);

Signal ProductNode_Float131Output_162: float (5 downto -14);
Signal ProductNode_Float132weight : float ( 5 downto -14 ) := to_float (0.985013,5,14);

Signal ProductNode_Float132Output_163: float (5 downto -14);
Signal ProductNode_Float133weight : float ( 5 downto -14 ) := to_float (0.592017,5,14);

Signal ProductNode_Float133Output_164: float (5 downto -14);
Signal SumNode_Float31Output_165: float (5 downto -14);
Signal ProductNode_Float134Output_166: float (5 downto -14);
Signal SumNode_Float32Output_167: float (5 downto -14);
Signal ProductNode_Float135Output_168: float (5 downto -14);
Signal ProductNode_Float136weight : float ( 5 downto -14 ) := to_float (0.479802,5,14);

Signal ProductNode_Float136Output_169: float (5 downto -14);
Signal SumNode_Float33Output_170: float (5 downto -14);
Signal ProductNode_Float137Output_171: float (5 downto -14);
Signal ProductNode_Float138weight : float ( 5 downto -14 ) := to_float (0.927615,5,14);

Signal ProductNode_Float138Output_172: float (5 downto -14);
Signal ProductNode_Float139weight : float ( 5 downto -14 ) := to_float (0.792795,5,14);

Signal ProductNode_Float139Output_173: float (5 downto -14);
Signal SumNode_Float34Output_174: float (5 downto -14);
Signal ProductNode_Float140Output_175: float (5 downto -14);
Signal ProductNode_Float141weight : float ( 5 downto -14 ) := to_float (0.907425,5,14);

Signal ProductNode_Float141Output_176: float (5 downto -14);
Signal ProductNode_Float142weight : float ( 5 downto -14 ) := to_float (0.948402,5,14);

Signal ProductNode_Float142Output_177: float (5 downto -14);
Signal ProductNode_Float143weight : float ( 5 downto -14 ) := to_float (0.838940,5,14);

Signal ProductNode_Float143Output_178: float (5 downto -14);
Signal ProductNode_Float144weight : float ( 5 downto -14 ) := to_float (0.898142,5,14);

Signal ProductNode_Float144Output_179: float (5 downto -14);
Signal SumNode_Float35Output_180: float (5 downto -14);
Signal ProductNode_Float145Output_181: float (5 downto -14);
Signal ProductNode_Float146weight : float ( 5 downto -14 ) := to_float (0.826105,5,14);

Signal ProductNode_Float146Output_182: float (5 downto -14);
Signal ProductNode_Float147weight : float ( 5 downto -14 ) := to_float (0.838083,5,14);

Signal ProductNode_Float147Output_183: float (5 downto -14);
Signal SumNode_Float36Output_184: float (5 downto -14);
Signal ProductNode_Float148Output_185: float (5 downto -14);
Signal ProductNode_Float149weight : float ( 5 downto -14 ) := to_float (0.970921,5,14);

Signal ProductNode_Float149Output_186: float (5 downto -14);
Signal ProductNode_Float150weight : float ( 5 downto -14 ) := to_float (0.672140,5,14);

Signal ProductNode_Float150Output_187: float (5 downto -14);
Signal SumNode_Float37Output_188: float (5 downto -14);
Signal ProductNode_Float151Output_189: float (5 downto -14);
Signal ProductNode_Float152weight : float ( 5 downto -14 ) := to_float (0.989270,5,14);

Signal ProductNode_Float152Output_190: float (5 downto -14);
Signal ProductNode_Float153weight : float ( 5 downto -14 ) := to_float (0.997554,5,14);

Signal ProductNode_Float153Output_191: float (5 downto -14);
Signal ProductNode_Float154weight : float ( 5 downto -14 ) := to_float (0.414069,5,14);

Signal ProductNode_Float154Output_192: float (5 downto -14);
Signal SumNode_Float38Output_193: float (5 downto -14);
Signal ProductNode_Float155Output_194: float (5 downto -14);
Signal ProductNode_Float156weight : float ( 5 downto -14 ) := to_float (0.853307,5,14);

Signal ProductNode_Float156Output_195: float (5 downto -14);
Signal ProductNode_Float157weight : float ( 5 downto -14 ) := to_float (0.886527,5,14);

Signal ProductNode_Float157Output_196: float (5 downto -14);
Signal SumNode_Float39Output_197: float (5 downto -14);
Signal ProductNode_Float158Output_198: float (5 downto -14);
Signal ProductNode_Float159weight : float ( 5 downto -14 ) := to_float (0.554692,5,14);

Signal ProductNode_Float159Output_199: float (5 downto -14);
Signal ProductNode_Float160weight : float ( 5 downto -14 ) := to_float (0.989739,5,14);

Signal ProductNode_Float160Output_200: float (5 downto -14);
Signal ProductNode_Float161weight : float ( 5 downto -14 ) := to_float (0.549861,5,14);

Signal ProductNode_Float161Output_201: float (5 downto -14);
Signal SumNode_Float40Output_202: float (5 downto -14);
Signal ProductNode_Float162Output_203: float (5 downto -14);
Signal SumNode_Float41Output_204: float (5 downto -14);
Signal ProductNode_Float163Output_205: float (5 downto -14);
Signal ProductNode_Float164weight : float ( 5 downto -14 ) := to_float (0.970629,5,14);

Signal ProductNode_Float164Output_206: float (5 downto -14);
Signal ProductNode_Float165weight : float ( 5 downto -14 ) := to_float (0.817897,5,14);

Signal ProductNode_Float165Output_207: float (5 downto -14);
Signal ProductNode_Float166weight : float ( 5 downto -14 ) := to_float (0.912886,5,14);

Signal ProductNode_Float166Output_208: float (5 downto -14);
Signal SumNode_Float42Output_209: float (5 downto -14);
Signal ProductNode_Float167Output_210: float (5 downto -14);
Signal ProductNode_Float168weight : float ( 5 downto -14 ) := to_float (0.976301,5,14);

Signal ProductNode_Float168Output_211: float (5 downto -14);
Signal ProductNode_Float169weight : float ( 5 downto -14 ) := to_float (0.988880,5,14);

Signal ProductNode_Float169Output_212: float (5 downto -14);
Signal ProductNode_Float170weight : float ( 5 downto -14 ) := to_float (0.558577,5,14);

Signal ProductNode_Float170Output_213: float (5 downto -14);
Signal SumNode_Float43Output_214: float (5 downto -14);
Signal ProductNode_Float171Output_215: float (5 downto -14);
Signal ProductNode_Float172weight : float ( 5 downto -14 ) := to_float (0.731617,5,14);

Signal ProductNode_Float172Output_216: float (5 downto -14);
Signal ProductNode_Float173weight : float ( 5 downto -14 ) := to_float (0.954043,5,14);

Signal ProductNode_Float173Output_217: float (5 downto -14);
Signal SumNode_Float44Output_218: float (5 downto -14);
Signal ProductNode_Float174Output_219: float (5 downto -14);
Signal ProductNode_Float175weight : float ( 5 downto -14 ) := to_float (0.646579,5,14);

Signal ProductNode_Float175Output_220: float (5 downto -14);
Signal ProductNode_Float176weight : float ( 5 downto -14 ) := to_float (0.985013,5,14);

Signal ProductNode_Float176Output_221: float (5 downto -14);
Signal ProductNode_Float177weight : float ( 5 downto -14 ) := to_float (0.592017,5,14);

Signal ProductNode_Float177Output_222: float (5 downto -14);
Signal SumNode_Float45Output_223: float (5 downto -14);
Signal ProductNode_Float178Output_224: float (5 downto -14);
Signal SumNode_Float46Output_225: float (5 downto -14);
Signal ProductNode_Float179Output_226: float (5 downto -14);
Signal ProductNode_Float180weight : float ( 5 downto -14 ) := to_float (0.673404,5,14);

Signal ProductNode_Float180Output_227: float (5 downto -14);
Signal SumNode_Float47Output_228: float (5 downto -14);
Signal ProductNode_Float181Output_229: float (5 downto -14);
Signal ProductNode_Float182weight : float ( 5 downto -14 ) := to_float (0.750079,5,14);

Signal ProductNode_Float182Output_230: float (5 downto -14);
Signal ProductNode_Float183weight : float ( 5 downto -14 ) := to_float (0.947231,5,14);

Signal ProductNode_Float183Output_231: float (5 downto -14);
Signal SumNode_Float48Output_232: float (5 downto -14);
Signal ProductNode_Float184Output_233: float (5 downto -14);
Signal ProductNode_Float185weight : float ( 5 downto -14 ) := to_float (0.907425,5,14);

Signal ProductNode_Float185Output_234: float (5 downto -14);
Signal ProductNode_Float186weight : float ( 5 downto -14 ) := to_float (0.747070,5,14);

Signal ProductNode_Float186Output_235: float (5 downto -14);
Signal ProductNode_Float187weight : float ( 5 downto -14 ) := to_float (0.617466,5,14);

Signal ProductNode_Float187Output_236: float (5 downto -14);
Signal ProductNode_Float188weight : float ( 5 downto -14 ) := to_float (0.981367,5,14);

Signal ProductNode_Float188Output_237: float (5 downto -14);
Signal SumNode_Float49Output_238: float (5 downto -14);
Signal ProductNode_Float189Output_239: float (5 downto -14);
Signal ProductNode_Float190weight : float ( 5 downto -14 ) := to_float (0.826105,5,14);

Signal ProductNode_Float190Output_240: float (5 downto -14);
Signal ProductNode_Float191weight : float ( 5 downto -14 ) := to_float (0.898792,5,14);

Signal ProductNode_Float191Output_241: float (5 downto -14);
Signal SumNode_Float50Output_242: float (5 downto -14);
Signal ProductNode_Float192Output_243: float (5 downto -14);
Signal SumNode_Float51Output_244: float (5 downto -14);
Signal ProductNode_Float193Output_245: float (5 downto -14);
Signal ProductNode_Float194weight : float ( 5 downto -14 ) := to_float (0.995408,5,14);

Signal ProductNode_Float194Output_246: float (5 downto -14);
Signal ProductNode_Float195weight : float ( 5 downto -14 ) := to_float (0.970921,5,14);

Signal ProductNode_Float195Output_247: float (5 downto -14);
Signal ProductNode_Float196weight : float ( 5 downto -14 ) := to_float (0.672140,5,14);

Signal ProductNode_Float196Output_248: float (5 downto -14);
Signal SumNode_Float52Output_249: float (5 downto -14);
Signal ProductNode_Float197Output_250: float (5 downto -14);
Signal ProductNode_Float198weight : float ( 5 downto -14 ) := to_float (0.989270,5,14);

Signal ProductNode_Float198Output_251: float (5 downto -14);
Signal ProductNode_Float199weight : float ( 5 downto -14 ) := to_float (0.966381,5,14);

Signal ProductNode_Float199Output_252: float (5 downto -14);
Signal ProductNode_Float200weight : float ( 5 downto -14 ) := to_float (0.690672,5,14);

Signal ProductNode_Float200Output_253: float (5 downto -14);
Signal SumNode_Float53Output_254: float (5 downto -14);
Signal ProductNode_Float201Output_255: float (5 downto -14);
Signal ProductNode_Float202weight : float ( 5 downto -14 ) := to_float (0.853307,5,14);

Signal ProductNode_Float202Output_256: float (5 downto -14);
Signal ProductNode_Float203weight : float ( 5 downto -14 ) := to_float (0.886527,5,14);

Signal ProductNode_Float203Output_257: float (5 downto -14);
Signal SumNode_Float54Output_258: float (5 downto -14);
Signal ProductNode_Float204Output_259: float (5 downto -14);
Signal ProductNode_Float205weight : float ( 5 downto -14 ) := to_float (0.554692,5,14);

Signal ProductNode_Float205Output_260: float (5 downto -14);
Signal ProductNode_Float206weight : float ( 5 downto -14 ) := to_float (0.941870,5,14);

Signal ProductNode_Float206Output_261: float (5 downto -14);
Signal ProductNode_Float207weight : float ( 5 downto -14 ) := to_float (0.763101,5,14);

Signal ProductNode_Float207Output_262: float (5 downto -14);
Signal SumNode_Float55Output_263: float (5 downto -14);
Signal ProductNode_Float208Output_264: float (5 downto -14);
Signal SumNode_Float56Output_265: float (5 downto -14);
Signal ProductNode_Float209Output_266: float (5 downto -14);
Signal ProductNode_Float210weight : float ( 5 downto -14 ) := to_float (0.951966,5,14);

Signal ProductNode_Float210Output_267: float (5 downto -14);
Signal ProductNode_Float211weight : float ( 5 downto -14 ) := to_float (0.817897,5,14);

Signal ProductNode_Float211Output_268: float (5 downto -14);
Signal ProductNode_Float212weight : float ( 5 downto -14 ) := to_float (0.912886,5,14);

Signal ProductNode_Float212Output_269: float (5 downto -14);
Signal SumNode_Float57Output_270: float (5 downto -14);
Signal ProductNode_Float213Output_271: float (5 downto -14);
Signal ProductNode_Float214weight : float ( 5 downto -14 ) := to_float (0.976301,5,14);

Signal ProductNode_Float214Output_272: float (5 downto -14);
Signal ProductNode_Float215weight : float ( 5 downto -14 ) := to_float (0.909585,5,14);

Signal ProductNode_Float215Output_273: float (5 downto -14);
Signal ProductNode_Float216weight : float ( 5 downto -14 ) := to_float (0.822920,5,14);

Signal ProductNode_Float216Output_274: float (5 downto -14);
Signal SumNode_Float58Output_275: float (5 downto -14);
Signal ProductNode_Float217Output_276: float (5 downto -14);
Signal ProductNode_Float218weight : float ( 5 downto -14 ) := to_float (0.731617,5,14);

Signal ProductNode_Float218Output_277: float (5 downto -14);
Signal ProductNode_Float219weight : float ( 5 downto -14 ) := to_float (0.954043,5,14);

Signal ProductNode_Float219Output_278: float (5 downto -14);
Signal SumNode_Float59Output_279: float (5 downto -14);
Signal ProductNode_Float220Output_280: float (5 downto -14);
Signal ProductNode_Float221weight : float ( 5 downto -14 ) := to_float (0.646579,5,14);

Signal ProductNode_Float221Output_281: float (5 downto -14);
Signal ProductNode_Float222weight : float ( 5 downto -14 ) := to_float (0.790147,5,14);

Signal ProductNode_Float222Output_282: float (5 downto -14);
Signal ProductNode_Float223weight : float ( 5 downto -14 ) := to_float (0.929014,5,14);

Signal ProductNode_Float223Output_283: float (5 downto -14);
Signal SumNode_Float60Output_284: float (5 downto -14);
Signal ProductNode_Float224Output_285: float (5 downto -14);
Signal SumNode_Float61Output_286: float (5 downto -14);
Signal ProductNode_Float225Output_287: float (5 downto -14);
Signal ProductNode_Float226weight : float ( 5 downto -14 ) := to_float (0.737500,5,14);

Signal ProductNode_Float226Output_288: float (5 downto -14);
Signal SumNode_Float62Output_289: float (5 downto -14);
Signal ProductNode_Float227Output_290: float (5 downto -14);
Signal ProductNode_Float228weight : float ( 5 downto -14 ) := to_float (0.927615,5,14);

Signal ProductNode_Float228Output_291: float (5 downto -14);
Signal ProductNode_Float229weight : float ( 5 downto -14 ) := to_float (0.792795,5,14);

Signal ProductNode_Float229Output_292: float (5 downto -14);
Signal SumNode_Float63Output_293: float (5 downto -14);
Signal ProductNode_Float230Output_294: float (5 downto -14);
Signal ProductNode_Float231weight : float ( 5 downto -14 ) := to_float (0.807766,5,14);

Signal ProductNode_Float231Output_295: float (5 downto -14);
Signal ProductNode_Float232weight : float ( 5 downto -14 ) := to_float (0.907576,5,14);

Signal ProductNode_Float232Output_296: float (5 downto -14);
Signal ProductNode_Float233weight : float ( 5 downto -14 ) := to_float (0.838940,5,14);

Signal ProductNode_Float233Output_297: float (5 downto -14);
Signal ProductNode_Float234weight : float ( 5 downto -14 ) := to_float (0.898142,5,14);

Signal ProductNode_Float234Output_298: float (5 downto -14);
Signal SumNode_Float64Output_299: float (5 downto -14);
Signal ProductNode_Float235Output_300: float (5 downto -14);
Signal ProductNode_Float236weight : float ( 5 downto -14 ) := to_float (0.919167,5,14);

Signal ProductNode_Float236Output_301: float (5 downto -14);
Signal ProductNode_Float237weight : float ( 5 downto -14 ) := to_float (0.781132,5,14);

Signal ProductNode_Float237Output_302: float (5 downto -14);
Signal SumNode_Float65Output_303: float (5 downto -14);
Signal ProductNode_Float238Output_304: float (5 downto -14);
Signal ProductNode_Float239weight : float ( 5 downto -14 ) := to_float (0.970921,5,14);

Signal ProductNode_Float239Output_305: float (5 downto -14);
Signal ProductNode_Float240weight : float ( 5 downto -14 ) := to_float (0.672140,5,14);

Signal ProductNode_Float240Output_306: float (5 downto -14);
Signal SumNode_Float66Output_307: float (5 downto -14);
Signal ProductNode_Float241Output_308: float (5 downto -14);
Signal ProductNode_Float242weight : float ( 5 downto -14 ) := to_float (0.989270,5,14);

Signal ProductNode_Float242Output_309: float (5 downto -14);
Signal ProductNode_Float243weight : float ( 5 downto -14 ) := to_float (0.966381,5,14);

Signal ProductNode_Float243Output_310: float (5 downto -14);
Signal ProductNode_Float244weight : float ( 5 downto -14 ) := to_float (0.690672,5,14);

Signal ProductNode_Float244Output_311: float (5 downto -14);
Signal SumNode_Float67Output_312: float (5 downto -14);
Signal ProductNode_Float245Output_313: float (5 downto -14);
Signal ProductNode_Float246weight : float ( 5 downto -14 ) := to_float (0.853307,5,14);

Signal ProductNode_Float246Output_314: float (5 downto -14);
Signal ProductNode_Float247weight : float ( 5 downto -14 ) := to_float (0.886527,5,14);

Signal ProductNode_Float247Output_315: float (5 downto -14);
Signal SumNode_Float68Output_316: float (5 downto -14);
Signal ProductNode_Float248Output_317: float (5 downto -14);
Signal ProductNode_Float249weight : float ( 5 downto -14 ) := to_float (0.554692,5,14);

Signal ProductNode_Float249Output_318: float (5 downto -14);
Signal ProductNode_Float250weight : float ( 5 downto -14 ) := to_float (0.941870,5,14);

Signal ProductNode_Float250Output_319: float (5 downto -14);
Signal ProductNode_Float251weight : float ( 5 downto -14 ) := to_float (0.763101,5,14);

Signal ProductNode_Float251Output_320: float (5 downto -14);
Signal SumNode_Float69Output_321: float (5 downto -14);
Signal ProductNode_Float252Output_322: float (5 downto -14);
Signal SumNode_Float70Output_323: float (5 downto -14);
Signal ProductNode_Float253Output_324: float (5 downto -14);
Signal ProductNode_Float254weight : float ( 5 downto -14 ) := to_float (0.840616,5,14);

Signal ProductNode_Float254Output_325: float (5 downto -14);
Signal ProductNode_Float255weight : float ( 5 downto -14 ) := to_float (0.817897,5,14);

Signal ProductNode_Float255Output_326: float (5 downto -14);
Signal ProductNode_Float256weight : float ( 5 downto -14 ) := to_float (0.912886,5,14);

Signal ProductNode_Float256Output_327: float (5 downto -14);
Signal SumNode_Float71Output_328: float (5 downto -14);
Signal ProductNode_Float257Output_329: float (5 downto -14);
Signal ProductNode_Float258weight : float ( 5 downto -14 ) := to_float (0.976301,5,14);

Signal ProductNode_Float258Output_330: float (5 downto -14);
Signal ProductNode_Float259weight : float ( 5 downto -14 ) := to_float (0.909585,5,14);

Signal ProductNode_Float259Output_331: float (5 downto -14);
Signal ProductNode_Float260weight : float ( 5 downto -14 ) := to_float (0.822920,5,14);

Signal ProductNode_Float260Output_332: float (5 downto -14);
Signal SumNode_Float72Output_333: float (5 downto -14);
Signal ProductNode_Float261Output_334: float (5 downto -14);
Signal ProductNode_Float262weight : float ( 5 downto -14 ) := to_float (0.731617,5,14);

Signal ProductNode_Float262Output_335: float (5 downto -14);
Signal ProductNode_Float263weight : float ( 5 downto -14 ) := to_float (0.954043,5,14);

Signal ProductNode_Float263Output_336: float (5 downto -14);
Signal SumNode_Float73Output_337: float (5 downto -14);
Signal ProductNode_Float264Output_338: float (5 downto -14);
Signal ProductNode_Float265weight : float ( 5 downto -14 ) := to_float (0.646579,5,14);

Signal ProductNode_Float265Output_339: float (5 downto -14);
Signal ProductNode_Float266weight : float ( 5 downto -14 ) := to_float (0.790147,5,14);

Signal ProductNode_Float266Output_340: float (5 downto -14);
Signal ProductNode_Float267weight : float ( 5 downto -14 ) := to_float (0.929014,5,14);

Signal ProductNode_Float267Output_341: float (5 downto -14);
Signal SumNode_Float74Output_342: float (5 downto -14);
Signal ProductNode_Float268Output_343: float (5 downto -14);
Signal SumNode_Float75Output_344: float (5 downto -14);
Signal ProductNode_Float269Output_345: float (5 downto -14);
Signal ProductNode_Float270weight : float ( 5 downto -14 ) := to_float (0.896858,5,14);

Signal ProductNode_Float270Output_346: float (5 downto -14);
Signal SumNode_Float76Output_347: float (5 downto -14);
Signal ProductNode_Float271Output_348: float (5 downto -14);
Signal ProductNode_Float272weight : float ( 5 downto -14 ) := to_float (0.750079,5,14);

Signal ProductNode_Float272Output_349: float (5 downto -14);
Signal ProductNode_Float273weight : float ( 5 downto -14 ) := to_float (0.947231,5,14);

Signal ProductNode_Float273Output_350: float (5 downto -14);
Signal SumNode_Float77Output_351: float (5 downto -14);
Signal ProductNode_Float274Output_352: float (5 downto -14);
Signal ProductNode_Float275weight : float ( 5 downto -14 ) := to_float (0.807766,5,14);

Signal ProductNode_Float275Output_353: float (5 downto -14);
Signal ProductNode_Float276weight : float ( 5 downto -14 ) := to_float (0.825885,5,14);

Signal ProductNode_Float276Output_354: float (5 downto -14);
Signal ProductNode_Float277weight : float ( 5 downto -14 ) := to_float (0.617466,5,14);

Signal ProductNode_Float277Output_355: float (5 downto -14);
Signal ProductNode_Float278weight : float ( 5 downto -14 ) := to_float (0.981367,5,14);

Signal ProductNode_Float278Output_356: float (5 downto -14);
Signal SumNode_Float78Output_357: float (5 downto -14);
Signal ProductNode_Float279Output_358: float (5 downto -14);
Signal ProductNode_Float280weight : float ( 5 downto -14 ) := to_float (0.919167,5,14);

Signal ProductNode_Float280Output_359: float (5 downto -14);
Signal ProductNode_Float281weight : float ( 5 downto -14 ) := to_float (0.933580,5,14);

Signal ProductNode_Float281Output_360: float (5 downto -14);
Signal SumNode_Float79Output_361: float (5 downto -14);
Signal ProductNode_Float282Output_362: float (5 downto -14);
Signal SumNode_Float80Output_363: float (5 downto -14);
Signal ProductNode_Float283Output_364: float (5 downto -14);
Signal ProductNode_Float284weight : float ( 5 downto -14 ) := to_float (0.469245,5,14);

Signal ProductNode_Float284Output_365: float (5 downto -14);
Signal SumNode_Float81Output_366: float (5 downto -14);
Signal ProductNode_Float285Output_367: float (5 downto -14);
Signal ProductNode_Float286weight : float ( 5 downto -14 ) := to_float (0.848299,5,14);

Signal ProductNode_Float286Output_368: float (5 downto -14);
Signal ProductNode_Float287weight : float ( 5 downto -14 ) := to_float (0.895308,5,14);

Signal ProductNode_Float287Output_369: float (5 downto -14);
Signal ProductNode_Float288weight : float ( 5 downto -14 ) := to_float (0.842608,5,14);

Signal ProductNode_Float288Output_370: float (5 downto -14);
Signal SumNode_Float82Output_371: float (5 downto -14);
Signal ProductNode_Float289Output_372: float (5 downto -14);
Signal ProductNode_Float290weight : float ( 5 downto -14 ) := to_float (0.870697,5,14);

Signal ProductNode_Float290Output_373: float (5 downto -14);
Signal ProductNode_Float291weight : float ( 5 downto -14 ) := to_float (0.945793,5,14);

Signal ProductNode_Float291Output_374: float (5 downto -14);
Signal ProductNode_Float292weight : float ( 5 downto -14 ) := to_float (0.954870,5,14);

Signal ProductNode_Float292Output_375: float (5 downto -14);
Signal ProductNode_Float293weight : float ( 5 downto -14 ) := to_float (0.870404,5,14);

Signal ProductNode_Float293Output_376: float (5 downto -14);
Signal ProductNode_Float294weight : float ( 5 downto -14 ) := to_float (0.780732,5,14);

Signal ProductNode_Float294Output_377: float (5 downto -14);
Signal ProductNode_Float295weight : float ( 5 downto -14 ) := to_float (0.810846,5,14);

Signal ProductNode_Float295Output_378: float (5 downto -14);
Signal SumNode_Float83Output_379: float (5 downto -14);
Signal ProductNode_Float296Output_380: float (5 downto -14);
Signal ProductNode_Float297weight : float ( 5 downto -14 ) := to_float (0.991361,5,14);

Signal ProductNode_Float297Output_381: float (5 downto -14);
Signal ProductNode_Float298weight : float ( 5 downto -14 ) := to_float (0.669241,5,14);

Signal ProductNode_Float298Output_382: float (5 downto -14);
Signal ProductNode_Float299weight : float ( 5 downto -14 ) := to_float (0.971580,5,14);

Signal ProductNode_Float299Output_383: float (5 downto -14);
Signal SumNode_Float84Output_384: float (5 downto -14);
Signal ProductNode_Float300Output_385: float (5 downto -14);
Signal ProductNode_Float301weight : float ( 5 downto -14 ) := to_float (0.870697,5,14);

Signal ProductNode_Float301Output_386: float (5 downto -14);
Signal ProductNode_Float302weight : float ( 5 downto -14 ) := to_float (0.753690,5,14);

Signal ProductNode_Float302Output_387: float (5 downto -14);
Signal ProductNode_Float303weight : float ( 5 downto -14 ) := to_float (0.774480,5,14);

Signal ProductNode_Float303Output_388: float (5 downto -14);
Signal ProductNode_Float304weight : float ( 5 downto -14 ) := to_float (0.870404,5,14);

Signal ProductNode_Float304Output_389: float (5 downto -14);
Signal ProductNode_Float305weight : float ( 5 downto -14 ) := to_float (0.933776,5,14);

Signal ProductNode_Float305Output_390: float (5 downto -14);
Signal ProductNode_Float306weight : float ( 5 downto -14 ) := to_float (0.660973,5,14);

Signal ProductNode_Float306Output_391: float (5 downto -14);
Signal SumNode_Float85Output_392: float (5 downto -14);
Signal ProductNode_Float307Output_393: float (5 downto -14);
Signal ProductNode_Float308weight : float ( 5 downto -14 ) := to_float (0.870239,5,14);

Signal ProductNode_Float308Output_394: float (5 downto -14);
Signal SumNode_Float86Output_395: float (5 downto -14);
Signal ProductNode_Float309Output_396: float (5 downto -14);
Signal ProductNode_Float310weight : float ( 5 downto -14 ) := to_float (0.756327,5,14);

Signal ProductNode_Float310Output_397: float (5 downto -14);
Signal ProductNode_Float311weight : float ( 5 downto -14 ) := to_float (0.890735,5,14);

Signal ProductNode_Float311Output_398: float (5 downto -14);
Signal ProductNode_Float312weight : float ( 5 downto -14 ) := to_float (0.689002,5,14);

Signal ProductNode_Float312Output_399: float (5 downto -14);
Signal ProductNode_Float313weight : float ( 5 downto -14 ) := to_float (0.966814,5,14);

Signal ProductNode_Float313Output_400: float (5 downto -14);
Signal SumNode_Float87Output_401: float (5 downto -14);
Signal ProductNode_Float314Output_402: float (5 downto -14);
Signal ProductNode_Float315weight : float ( 5 downto -14 ) := to_float (0.551341,5,14);

Signal ProductNode_Float315Output_403: float (5 downto -14);
Signal ProductNode_Float316weight : float ( 5 downto -14 ) := to_float (0.795357,5,14);

Signal ProductNode_Float316Output_404: float (5 downto -14);
Signal ProductNode_Float317weight : float ( 5 downto -14 ) := to_float (0.746308,5,14);

Signal ProductNode_Float317Output_405: float (5 downto -14);
Signal ProductNode_Float318weight : float ( 5 downto -14 ) := to_float (0.989597,5,14);

Signal ProductNode_Float318Output_406: float (5 downto -14);
Signal ProductNode_Float319weight : float ( 5 downto -14 ) := to_float (0.577708,5,14);

Signal ProductNode_Float319Output_407: float (5 downto -14);
Signal ProductNode_Float320weight : float ( 5 downto -14 ) := to_float (0.618274,5,14);

Signal ProductNode_Float320Output_408: float (5 downto -14);
Signal SumNode_Float88Output_409: float (5 downto -14);
Signal ProductNode_Float321Output_410: float (5 downto -14);
Signal ProductNode_Float322weight : float ( 5 downto -14 ) := to_float (0.952809,5,14);

Signal ProductNode_Float322Output_411: float (5 downto -14);
Signal ProductNode_Float323weight : float ( 5 downto -14 ) := to_float (0.495915,5,14);

Signal ProductNode_Float323Output_412: float (5 downto -14);
Signal ProductNode_Float324weight : float ( 5 downto -14 ) := to_float (0.993928,5,14);

Signal ProductNode_Float324Output_413: float (5 downto -14);
Signal SumNode_Float89Output_414: float (5 downto -14);
Signal ProductNode_Float325Output_415: float (5 downto -14);
Signal ProductNode_Float326weight : float ( 5 downto -14 ) := to_float (0.551341,5,14);

Signal ProductNode_Float326Output_416: float (5 downto -14);
Signal ProductNode_Float327weight : float ( 5 downto -14 ) := to_float (0.926235,5,14);

Signal ProductNode_Float327Output_417: float (5 downto -14);
Signal ProductNode_Float328weight : float ( 5 downto -14 ) := to_float (0.616494,5,14);

Signal ProductNode_Float328Output_418: float (5 downto -14);
Signal ProductNode_Float329weight : float ( 5 downto -14 ) := to_float (0.989597,5,14);

Signal ProductNode_Float329Output_419: float (5 downto -14);
Signal ProductNode_Float330weight : float ( 5 downto -14 ) := to_float (0.986786,5,14);

Signal ProductNode_Float330Output_420: float (5 downto -14);
Signal ProductNode_Float331weight : float ( 5 downto -14 ) := to_float (0.464416,5,14);

Signal ProductNode_Float331Output_421: float (5 downto -14);
Signal SumNode_Float90Output_422: float (5 downto -14);
Signal ProductNode_Float332Output_423: float (5 downto -14);
Signal ProductNode_Float333weight : float ( 5 downto -14 ) := to_float (0.770987,5,14);

Signal ProductNode_Float333Output_424: float (5 downto -14);
Signal SumNode_Float91Output_425: float (5 downto -14);
Signal ProductNode_Float334Output_426: float (5 downto -14);
Signal ProductNode_Float335weight : float ( 5 downto -14 ) := to_float (0.906302,5,14);

Signal ProductNode_Float335Output_427: float (5 downto -14);
Signal SumNode_Float92Output_428: float (5 downto -14);
Signal ProductNode_Float336Output_429: float (5 downto -14);
Signal ProductNode_Float337weight : float ( 5 downto -14 ) := to_float (0.800117,5,14);

Signal ProductNode_Float337Output_430: float (5 downto -14);
Signal ProductNode_Float338weight : float ( 5 downto -14 ) := to_float (0.848299,5,14);

Signal ProductNode_Float338Output_431: float (5 downto -14);
Signal ProductNode_Float339weight : float ( 5 downto -14 ) := to_float (0.562709,5,14);

Signal ProductNode_Float339Output_432: float (5 downto -14);
Signal ProductNode_Float340weight : float ( 5 downto -14 ) := to_float (0.988453,5,14);

Signal ProductNode_Float340Output_433: float (5 downto -14);
Signal SumNode_Float93Output_434: float (5 downto -14);
Signal ProductNode_Float341Output_435: float (5 downto -14);
Signal ProductNode_Float342weight : float ( 5 downto -14 ) := to_float (0.870697,5,14);

Signal ProductNode_Float342Output_436: float (5 downto -14);
Signal ProductNode_Float343weight : float ( 5 downto -14 ) := to_float (0.945793,5,14);

Signal ProductNode_Float343Output_437: float (5 downto -14);
Signal ProductNode_Float344weight : float ( 5 downto -14 ) := to_float (0.729204,5,14);

Signal ProductNode_Float344Output_438: float (5 downto -14);
Signal ProductNode_Float345weight : float ( 5 downto -14 ) := to_float (0.870404,5,14);

Signal ProductNode_Float345Output_439: float (5 downto -14);
Signal ProductNode_Float346weight : float ( 5 downto -14 ) := to_float (0.780732,5,14);

Signal ProductNode_Float346Output_440: float (5 downto -14);
Signal ProductNode_Float347weight : float ( 5 downto -14 ) := to_float (0.917308,5,14);

Signal ProductNode_Float347Output_441: float (5 downto -14);
Signal SumNode_Float94Output_442: float (5 downto -14);
Signal ProductNode_Float348Output_443: float (5 downto -14);
Signal ProductNode_Float349weight : float ( 5 downto -14 ) := to_float (0.979033,5,14);

Signal ProductNode_Float349Output_444: float (5 downto -14);
Signal ProductNode_Float350weight : float ( 5 downto -14 ) := to_float (0.453222,5,14);

Signal ProductNode_Float350Output_445: float (5 downto -14);
Signal ProductNode_Float351weight : float ( 5 downto -14 ) := to_float (0.996146,5,14);

Signal ProductNode_Float351Output_446: float (5 downto -14);
Signal SumNode_Float95Output_447: float (5 downto -14);
Signal ProductNode_Float352Output_448: float (5 downto -14);
Signal ProductNode_Float353weight : float ( 5 downto -14 ) := to_float (0.870697,5,14);

Signal ProductNode_Float353Output_449: float (5 downto -14);
Signal ProductNode_Float354weight : float ( 5 downto -14 ) := to_float (0.753690,5,14);

Signal ProductNode_Float354Output_450: float (5 downto -14);
Signal ProductNode_Float355weight : float ( 5 downto -14 ) := to_float (0.936763,5,14);

Signal ProductNode_Float355Output_451: float (5 downto -14);
Signal ProductNode_Float356weight : float ( 5 downto -14 ) := to_float (0.870404,5,14);

Signal ProductNode_Float356Output_452: float (5 downto -14);
Signal ProductNode_Float357weight : float ( 5 downto -14 ) := to_float (0.933776,5,14);

Signal ProductNode_Float357Output_453: float (5 downto -14);
Signal ProductNode_Float358weight : float ( 5 downto -14 ) := to_float (0.973389,5,14);

Signal ProductNode_Float358Output_454: float (5 downto -14);
Signal SumNode_Float96Output_455: float (5 downto -14);
Signal ProductNode_Float359Output_456: float (5 downto -14);
Signal ProductNode_Float360weight : float ( 5 downto -14 ) := to_float (0.818419,5,14);

Signal ProductNode_Float360Output_457: float (5 downto -14);
Signal SumNode_Float97Output_458: float (5 downto -14);
Signal ProductNode_Float361Output_459: float (5 downto -14);
Signal ProductNode_Float362weight : float ( 5 downto -14 ) := to_float (0.940496,5,14);

Signal ProductNode_Float362Output_460: float (5 downto -14);
Signal ProductNode_Float363weight : float ( 5 downto -14 ) := to_float (0.890735,5,14);

Signal ProductNode_Float363Output_461: float (5 downto -14);
Signal ProductNode_Float364weight : float ( 5 downto -14 ) := to_float (0.382644,5,14);

Signal ProductNode_Float364Output_462: float (5 downto -14);
Signal ProductNode_Float365weight : float ( 5 downto -14 ) := to_float (0.998354,5,14);

Signal ProductNode_Float365Output_463: float (5 downto -14);
Signal SumNode_Float98Output_464: float (5 downto -14);
Signal ProductNode_Float366Output_465: float (5 downto -14);
Signal ProductNode_Float367weight : float ( 5 downto -14 ) := to_float (0.551341,5,14);

Signal ProductNode_Float367Output_466: float (5 downto -14);
Signal ProductNode_Float368weight : float ( 5 downto -14 ) := to_float (0.795357,5,14);

Signal ProductNode_Float368Output_467: float (5 downto -14);
Signal ProductNode_Float369weight : float ( 5 downto -14 ) := to_float (0.948695,5,14);

Signal ProductNode_Float369Output_468: float (5 downto -14);
Signal ProductNode_Float370weight : float ( 5 downto -14 ) := to_float (0.989597,5,14);

Signal ProductNode_Float370Output_469: float (5 downto -14);
Signal ProductNode_Float371weight : float ( 5 downto -14 ) := to_float (0.577708,5,14);

Signal ProductNode_Float371Output_470: float (5 downto -14);
Signal ProductNode_Float372weight : float ( 5 downto -14 ) := to_float (0.981240,5,14);

Signal ProductNode_Float372Output_471: float (5 downto -14);
Signal SumNode_Float99Output_472: float (5 downto -14);
Signal ProductNode_Float373Output_473: float (5 downto -14);
Signal ProductNode_Float374weight : float ( 5 downto -14 ) := to_float (0.960334,5,14);

Signal ProductNode_Float374Output_474: float (5 downto -14);
Signal ProductNode_Float375weight : float ( 5 downto -14 ) := to_float (0.336149,5,14);

Signal ProductNode_Float375Output_475: float (5 downto -14);
Signal ProductNode_Float376weight : float ( 5 downto -14 ) := to_float (0.999140,5,14);

Signal ProductNode_Float376Output_476: float (5 downto -14);
Signal SumNode_Float100Output_477: float (5 downto -14);
Signal ProductNode_Float377Output_478: float (5 downto -14);
Signal ProductNode_Float378weight : float ( 5 downto -14 ) := to_float (0.551341,5,14);

Signal ProductNode_Float378Output_479: float (5 downto -14);
Signal ProductNode_Float379weight : float ( 5 downto -14 ) := to_float (0.926235,5,14);

Signal ProductNode_Float379Output_480: float (5 downto -14);
Signal ProductNode_Float380weight : float ( 5 downto -14 ) := to_float (0.981519,5,14);

Signal ProductNode_Float380Output_481: float (5 downto -14);
Signal ProductNode_Float381weight : float ( 5 downto -14 ) := to_float (0.989597,5,14);

Signal ProductNode_Float381Output_482: float (5 downto -14);
Signal ProductNode_Float382weight : float ( 5 downto -14 ) := to_float (0.986786,5,14);

Signal ProductNode_Float382Output_483: float (5 downto -14);
Signal ProductNode_Float383weight : float ( 5 downto -14 ) := to_float (0.995641,5,14);

Signal ProductNode_Float383Output_484: float (5 downto -14);
Signal SumNode_Float101Output_485: float (5 downto -14);
Signal ProductNode_Float384Output_486: float (5 downto -14);
Signal ProductNode_Float385weight : float ( 5 downto -14 ) := to_float (0.664315,5,14);

Signal ProductNode_Float385Output_487: float (5 downto -14);
Signal SumNode_Float102Output_488: float (5 downto -14);
Signal ProductNode_Float386Output_489: float (5 downto -14);
Signal ProductNode_Float387weight : float ( 5 downto -14 ) := to_float (0.978597,5,14);

Signal ProductNode_Float387Output_490: float (5 downto -14);
Signal SumNode_Float103Output_491: float (5 downto -14);
Signal ProductNode_Float388Output_492: float (5 downto -14);
Signal ProductNode_Float389weight : float ( 5 downto -14 ) := to_float (0.655866,5,14);

Signal ProductNode_Float389Output_493: float (5 downto -14);
Signal SumNode_Float104Output_494: float (5 downto -14);
Signal ProductNode_Float390Output_495: float (5 downto -14);
Signal ProductNode_Float391weight : float ( 5 downto -14 ) := to_float (0.970921,5,14);

Signal ProductNode_Float391Output_496: float (5 downto -14);
Signal ProductNode_Float392weight : float ( 5 downto -14 ) := to_float (0.672140,5,14);

Signal ProductNode_Float392Output_497: float (5 downto -14);
Signal SumNode_Float105Output_498: float (5 downto -14);
Signal ProductNode_Float393Output_499: float (5 downto -14);
Signal ProductNode_Float394weight : float ( 5 downto -14 ) := to_float (0.989270,5,14);

Signal ProductNode_Float394Output_500: float (5 downto -14);
Signal ProductNode_Float395weight : float ( 5 downto -14 ) := to_float (0.997554,5,14);

Signal ProductNode_Float395Output_501: float (5 downto -14);
Signal ProductNode_Float396weight : float ( 5 downto -14 ) := to_float (0.414069,5,14);

Signal ProductNode_Float396Output_502: float (5 downto -14);
Signal SumNode_Float106Output_503: float (5 downto -14);
Signal ProductNode_Float397Output_504: float (5 downto -14);
Signal ProductNode_Float398weight : float ( 5 downto -14 ) := to_float (0.853307,5,14);

Signal ProductNode_Float398Output_505: float (5 downto -14);
Signal ProductNode_Float399weight : float ( 5 downto -14 ) := to_float (0.886527,5,14);

Signal ProductNode_Float399Output_506: float (5 downto -14);
Signal SumNode_Float107Output_507: float (5 downto -14);
Signal ProductNode_Float400Output_508: float (5 downto -14);
Signal ProductNode_Float401weight : float ( 5 downto -14 ) := to_float (0.554692,5,14);

Signal ProductNode_Float401Output_509: float (5 downto -14);
Signal ProductNode_Float402weight : float ( 5 downto -14 ) := to_float (0.989739,5,14);

Signal ProductNode_Float402Output_510: float (5 downto -14);
Signal ProductNode_Float403weight : float ( 5 downto -14 ) := to_float (0.549861,5,14);

Signal ProductNode_Float403Output_511: float (5 downto -14);
Signal SumNode_Float108Output_512: float (5 downto -14);
Signal ProductNode_Float404Output_513: float (5 downto -14);
Signal SumNode_Float109Output_514: float (5 downto -14);
Signal ProductNode_Float405Output_515: float (5 downto -14);
Signal ProductNode_Float406weight : float ( 5 downto -14 ) := to_float (0.994862,5,14);

Signal ProductNode_Float406Output_516: float (5 downto -14);
Signal ProductNode_Float407weight : float ( 5 downto -14 ) := to_float (0.817897,5,14);

Signal ProductNode_Float407Output_517: float (5 downto -14);
Signal ProductNode_Float408weight : float ( 5 downto -14 ) := to_float (0.912886,5,14);

Signal ProductNode_Float408Output_518: float (5 downto -14);
Signal SumNode_Float110Output_519: float (5 downto -14);
Signal ProductNode_Float409Output_520: float (5 downto -14);
Signal ProductNode_Float410weight : float ( 5 downto -14 ) := to_float (0.976301,5,14);

Signal ProductNode_Float410Output_521: float (5 downto -14);
Signal ProductNode_Float411weight : float ( 5 downto -14 ) := to_float (0.988880,5,14);

Signal ProductNode_Float411Output_522: float (5 downto -14);
Signal ProductNode_Float412weight : float ( 5 downto -14 ) := to_float (0.558577,5,14);

Signal ProductNode_Float412Output_523: float (5 downto -14);
Signal SumNode_Float111Output_524: float (5 downto -14);
Signal ProductNode_Float413Output_525: float (5 downto -14);
Signal ProductNode_Float414weight : float ( 5 downto -14 ) := to_float (0.731617,5,14);

Signal ProductNode_Float414Output_526: float (5 downto -14);
Signal ProductNode_Float415weight : float ( 5 downto -14 ) := to_float (0.954043,5,14);

Signal ProductNode_Float415Output_527: float (5 downto -14);
Signal SumNode_Float112Output_528: float (5 downto -14);
Signal ProductNode_Float416Output_529: float (5 downto -14);
Signal ProductNode_Float417weight : float ( 5 downto -14 ) := to_float (0.646579,5,14);

Signal ProductNode_Float417Output_530: float (5 downto -14);
Signal ProductNode_Float418weight : float ( 5 downto -14 ) := to_float (0.985013,5,14);

Signal ProductNode_Float418Output_531: float (5 downto -14);
Signal ProductNode_Float419weight : float ( 5 downto -14 ) := to_float (0.592017,5,14);

Signal ProductNode_Float419Output_532: float (5 downto -14);
Signal SumNode_Float113Output_533: float (5 downto -14);
Signal ProductNode_Float420Output_534: float (5 downto -14);
Signal SumNode_Float114Output_535: float (5 downto -14);
Signal ProductNode_Float421Output_536: float (5 downto -14);
Signal ProductNode_Float422weight : float ( 5 downto -14 ) := to_float (0.479802,5,14);

Signal ProductNode_Float422Output_537: float (5 downto -14);
Signal SumNode_Float115Output_538: float (5 downto -14);
Signal ProductNode_Float423Output_539: float (5 downto -14);
Signal ProductNode_Float424weight : float ( 5 downto -14 ) := to_float (0.927615,5,14);

Signal ProductNode_Float424Output_540: float (5 downto -14);
Signal ProductNode_Float425weight : float ( 5 downto -14 ) := to_float (0.792795,5,14);

Signal ProductNode_Float425Output_541: float (5 downto -14);
Signal SumNode_Float116Output_542: float (5 downto -14);
Signal ProductNode_Float426Output_543: float (5 downto -14);
Signal ProductNode_Float427weight : float ( 5 downto -14 ) := to_float (0.907425,5,14);

Signal ProductNode_Float427Output_544: float (5 downto -14);
Signal ProductNode_Float428weight : float ( 5 downto -14 ) := to_float (0.948402,5,14);

Signal ProductNode_Float428Output_545: float (5 downto -14);
Signal ProductNode_Float429weight : float ( 5 downto -14 ) := to_float (0.838940,5,14);

Signal ProductNode_Float429Output_546: float (5 downto -14);
Signal ProductNode_Float430weight : float ( 5 downto -14 ) := to_float (0.898142,5,14);

Signal ProductNode_Float430Output_547: float (5 downto -14);
Signal SumNode_Float117Output_548: float (5 downto -14);
Signal ProductNode_Float431Output_549: float (5 downto -14);
Signal ProductNode_Float432weight : float ( 5 downto -14 ) := to_float (0.826105,5,14);

Signal ProductNode_Float432Output_550: float (5 downto -14);
Signal ProductNode_Float433weight : float ( 5 downto -14 ) := to_float (0.838083,5,14);

Signal ProductNode_Float433Output_551: float (5 downto -14);
Signal SumNode_Float118Output_552: float (5 downto -14);
Signal ProductNode_Float434Output_553: float (5 downto -14);
Signal ProductNode_Float435weight : float ( 5 downto -14 ) := to_float (0.970921,5,14);

Signal ProductNode_Float435Output_554: float (5 downto -14);
Signal ProductNode_Float436weight : float ( 5 downto -14 ) := to_float (0.672140,5,14);

Signal ProductNode_Float436Output_555: float (5 downto -14);
Signal SumNode_Float119Output_556: float (5 downto -14);
Signal ProductNode_Float437Output_557: float (5 downto -14);
Signal ProductNode_Float438weight : float ( 5 downto -14 ) := to_float (0.989270,5,14);

Signal ProductNode_Float438Output_558: float (5 downto -14);
Signal ProductNode_Float439weight : float ( 5 downto -14 ) := to_float (0.997554,5,14);

Signal ProductNode_Float439Output_559: float (5 downto -14);
Signal ProductNode_Float440weight : float ( 5 downto -14 ) := to_float (0.414069,5,14);

Signal ProductNode_Float440Output_560: float (5 downto -14);
Signal SumNode_Float120Output_561: float (5 downto -14);
Signal ProductNode_Float441Output_562: float (5 downto -14);
Signal ProductNode_Float442weight : float ( 5 downto -14 ) := to_float (0.853307,5,14);

Signal ProductNode_Float442Output_563: float (5 downto -14);
Signal ProductNode_Float443weight : float ( 5 downto -14 ) := to_float (0.886527,5,14);

Signal ProductNode_Float443Output_564: float (5 downto -14);
Signal SumNode_Float121Output_565: float (5 downto -14);
Signal ProductNode_Float444Output_566: float (5 downto -14);
Signal ProductNode_Float445weight : float ( 5 downto -14 ) := to_float (0.554692,5,14);

Signal ProductNode_Float445Output_567: float (5 downto -14);
Signal ProductNode_Float446weight : float ( 5 downto -14 ) := to_float (0.989739,5,14);

Signal ProductNode_Float446Output_568: float (5 downto -14);
Signal ProductNode_Float447weight : float ( 5 downto -14 ) := to_float (0.549861,5,14);

Signal ProductNode_Float447Output_569: float (5 downto -14);
Signal SumNode_Float122Output_570: float (5 downto -14);
Signal ProductNode_Float448Output_571: float (5 downto -14);
Signal SumNode_Float123Output_572: float (5 downto -14);
Signal ProductNode_Float449Output_573: float (5 downto -14);
Signal ProductNode_Float450weight : float ( 5 downto -14 ) := to_float (0.970629,5,14);

Signal ProductNode_Float450Output_574: float (5 downto -14);
Signal ProductNode_Float451weight : float ( 5 downto -14 ) := to_float (0.817897,5,14);

Signal ProductNode_Float451Output_575: float (5 downto -14);
Signal ProductNode_Float452weight : float ( 5 downto -14 ) := to_float (0.912886,5,14);

Signal ProductNode_Float452Output_576: float (5 downto -14);
Signal SumNode_Float124Output_577: float (5 downto -14);
Signal ProductNode_Float453Output_578: float (5 downto -14);
Signal ProductNode_Float454weight : float ( 5 downto -14 ) := to_float (0.976301,5,14);

Signal ProductNode_Float454Output_579: float (5 downto -14);
Signal ProductNode_Float455weight : float ( 5 downto -14 ) := to_float (0.988880,5,14);

Signal ProductNode_Float455Output_580: float (5 downto -14);
Signal ProductNode_Float456weight : float ( 5 downto -14 ) := to_float (0.558577,5,14);

Signal ProductNode_Float456Output_581: float (5 downto -14);
Signal SumNode_Float125Output_582: float (5 downto -14);
Signal ProductNode_Float457Output_583: float (5 downto -14);
Signal ProductNode_Float458weight : float ( 5 downto -14 ) := to_float (0.731617,5,14);

Signal ProductNode_Float458Output_584: float (5 downto -14);
Signal ProductNode_Float459weight : float ( 5 downto -14 ) := to_float (0.954043,5,14);

Signal ProductNode_Float459Output_585: float (5 downto -14);
Signal SumNode_Float126Output_586: float (5 downto -14);
Signal ProductNode_Float460Output_587: float (5 downto -14);
Signal ProductNode_Float461weight : float ( 5 downto -14 ) := to_float (0.646579,5,14);

Signal ProductNode_Float461Output_588: float (5 downto -14);
Signal ProductNode_Float462weight : float ( 5 downto -14 ) := to_float (0.985013,5,14);

Signal ProductNode_Float462Output_589: float (5 downto -14);
Signal ProductNode_Float463weight : float ( 5 downto -14 ) := to_float (0.592017,5,14);

Signal ProductNode_Float463Output_590: float (5 downto -14);
Signal SumNode_Float127Output_591: float (5 downto -14);
Signal ProductNode_Float464Output_592: float (5 downto -14);
Signal SumNode_Float128Output_593: float (5 downto -14);
Signal ProductNode_Float465Output_594: float (5 downto -14);
Signal ProductNode_Float466weight : float ( 5 downto -14 ) := to_float (0.673404,5,14);

Signal ProductNode_Float466Output_595: float (5 downto -14);
Signal SumNode_Float129Output_596: float (5 downto -14);
Signal ProductNode_Float467Output_597: float (5 downto -14);
Signal ProductNode_Float468weight : float ( 5 downto -14 ) := to_float (0.750079,5,14);

Signal ProductNode_Float468Output_598: float (5 downto -14);
Signal ProductNode_Float469weight : float ( 5 downto -14 ) := to_float (0.947231,5,14);

Signal ProductNode_Float469Output_599: float (5 downto -14);
Signal SumNode_Float130Output_600: float (5 downto -14);
Signal ProductNode_Float470Output_601: float (5 downto -14);
Signal ProductNode_Float471weight : float ( 5 downto -14 ) := to_float (0.907425,5,14);

Signal ProductNode_Float471Output_602: float (5 downto -14);
Signal ProductNode_Float472weight : float ( 5 downto -14 ) := to_float (0.747070,5,14);

Signal ProductNode_Float472Output_603: float (5 downto -14);
Signal ProductNode_Float473weight : float ( 5 downto -14 ) := to_float (0.617466,5,14);

Signal ProductNode_Float473Output_604: float (5 downto -14);
Signal ProductNode_Float474weight : float ( 5 downto -14 ) := to_float (0.981367,5,14);

Signal ProductNode_Float474Output_605: float (5 downto -14);
Signal SumNode_Float131Output_606: float (5 downto -14);
Signal ProductNode_Float475Output_607: float (5 downto -14);
Signal ProductNode_Float476weight : float ( 5 downto -14 ) := to_float (0.826105,5,14);

Signal ProductNode_Float476Output_608: float (5 downto -14);
Signal ProductNode_Float477weight : float ( 5 downto -14 ) := to_float (0.898792,5,14);

Signal ProductNode_Float477Output_609: float (5 downto -14);
Signal SumNode_Float132Output_610: float (5 downto -14);
Signal ProductNode_Float478Output_611: float (5 downto -14);
Signal SumNode_Float133Output_612: float (5 downto -14);
Signal ProductNode_Float479Output_613: float (5 downto -14);
Signal ProductNode_Float480weight : float ( 5 downto -14 ) := to_float (0.935776,5,14);

Signal ProductNode_Float480Output_614: float (5 downto -14);
Signal ProductNode_Float481weight : float ( 5 downto -14 ) := to_float (0.970921,5,14);

Signal ProductNode_Float481Output_615: float (5 downto -14);
Signal ProductNode_Float482weight : float ( 5 downto -14 ) := to_float (0.672140,5,14);

Signal ProductNode_Float482Output_616: float (5 downto -14);
Signal SumNode_Float134Output_617: float (5 downto -14);
Signal ProductNode_Float483Output_618: float (5 downto -14);
Signal ProductNode_Float484weight : float ( 5 downto -14 ) := to_float (0.989270,5,14);

Signal ProductNode_Float484Output_619: float (5 downto -14);
Signal ProductNode_Float485weight : float ( 5 downto -14 ) := to_float (0.966381,5,14);

Signal ProductNode_Float485Output_620: float (5 downto -14);
Signal ProductNode_Float486weight : float ( 5 downto -14 ) := to_float (0.690672,5,14);

Signal ProductNode_Float486Output_621: float (5 downto -14);
Signal SumNode_Float135Output_622: float (5 downto -14);
Signal ProductNode_Float487Output_623: float (5 downto -14);
Signal ProductNode_Float488weight : float ( 5 downto -14 ) := to_float (0.853307,5,14);

Signal ProductNode_Float488Output_624: float (5 downto -14);
Signal ProductNode_Float489weight : float ( 5 downto -14 ) := to_float (0.886527,5,14);

Signal ProductNode_Float489Output_625: float (5 downto -14);
Signal SumNode_Float136Output_626: float (5 downto -14);
Signal ProductNode_Float490Output_627: float (5 downto -14);
Signal ProductNode_Float491weight : float ( 5 downto -14 ) := to_float (0.554692,5,14);

Signal ProductNode_Float491Output_628: float (5 downto -14);
Signal ProductNode_Float492weight : float ( 5 downto -14 ) := to_float (0.941870,5,14);

Signal ProductNode_Float492Output_629: float (5 downto -14);
Signal ProductNode_Float493weight : float ( 5 downto -14 ) := to_float (0.763101,5,14);

Signal ProductNode_Float493Output_630: float (5 downto -14);
Signal SumNode_Float137Output_631: float (5 downto -14);
Signal ProductNode_Float494Output_632: float (5 downto -14);
Signal SumNode_Float138Output_633: float (5 downto -14);
Signal ProductNode_Float495Output_634: float (5 downto -14);
Signal ProductNode_Float496weight : float ( 5 downto -14 ) := to_float (0.951966,5,14);

Signal ProductNode_Float496Output_635: float (5 downto -14);
Signal ProductNode_Float497weight : float ( 5 downto -14 ) := to_float (0.817897,5,14);

Signal ProductNode_Float497Output_636: float (5 downto -14);
Signal ProductNode_Float498weight : float ( 5 downto -14 ) := to_float (0.912886,5,14);

Signal ProductNode_Float498Output_637: float (5 downto -14);
Signal SumNode_Float139Output_638: float (5 downto -14);
Signal ProductNode_Float499Output_639: float (5 downto -14);
Signal ProductNode_Float500weight : float ( 5 downto -14 ) := to_float (0.976301,5,14);

Signal ProductNode_Float500Output_640: float (5 downto -14);
Signal ProductNode_Float501weight : float ( 5 downto -14 ) := to_float (0.909585,5,14);

Signal ProductNode_Float501Output_641: float (5 downto -14);
Signal ProductNode_Float502weight : float ( 5 downto -14 ) := to_float (0.822920,5,14);

Signal ProductNode_Float502Output_642: float (5 downto -14);
Signal SumNode_Float140Output_643: float (5 downto -14);
Signal ProductNode_Float503Output_644: float (5 downto -14);
Signal ProductNode_Float504weight : float ( 5 downto -14 ) := to_float (0.731617,5,14);

Signal ProductNode_Float504Output_645: float (5 downto -14);
Signal ProductNode_Float505weight : float ( 5 downto -14 ) := to_float (0.954043,5,14);

Signal ProductNode_Float505Output_646: float (5 downto -14);
Signal SumNode_Float141Output_647: float (5 downto -14);
Signal ProductNode_Float506Output_648: float (5 downto -14);
Signal ProductNode_Float507weight : float ( 5 downto -14 ) := to_float (0.646579,5,14);

Signal ProductNode_Float507Output_649: float (5 downto -14);
Signal ProductNode_Float508weight : float ( 5 downto -14 ) := to_float (0.790147,5,14);

Signal ProductNode_Float508Output_650: float (5 downto -14);
Signal ProductNode_Float509weight : float ( 5 downto -14 ) := to_float (0.929014,5,14);

Signal ProductNode_Float509Output_651: float (5 downto -14);
Signal SumNode_Float142Output_652: float (5 downto -14);
Signal ProductNode_Float510Output_653: float (5 downto -14);
Signal SumNode_Float143Output_654: float (5 downto -14);
Signal ProductNode_Float511Output_655: float (5 downto -14);
Signal ProductNode_Float512weight : float ( 5 downto -14 ) := to_float (0.737500,5,14);

Signal ProductNode_Float512Output_656: float (5 downto -14);
Signal SumNode_Float144Output_657: float (5 downto -14);
Signal ProductNode_Float513Output_658: float (5 downto -14);
Signal ProductNode_Float514weight : float ( 5 downto -14 ) := to_float (0.927615,5,14);

Signal ProductNode_Float514Output_659: float (5 downto -14);
Signal ProductNode_Float515weight : float ( 5 downto -14 ) := to_float (0.792795,5,14);

Signal ProductNode_Float515Output_660: float (5 downto -14);
Signal SumNode_Float145Output_661: float (5 downto -14);
Signal ProductNode_Float516Output_662: float (5 downto -14);
Signal ProductNode_Float517weight : float ( 5 downto -14 ) := to_float (0.807766,5,14);

Signal ProductNode_Float517Output_663: float (5 downto -14);
Signal ProductNode_Float518weight : float ( 5 downto -14 ) := to_float (0.907576,5,14);

Signal ProductNode_Float518Output_664: float (5 downto -14);
Signal ProductNode_Float519weight : float ( 5 downto -14 ) := to_float (0.838940,5,14);

Signal ProductNode_Float519Output_665: float (5 downto -14);
Signal ProductNode_Float520weight : float ( 5 downto -14 ) := to_float (0.898142,5,14);

Signal ProductNode_Float520Output_666: float (5 downto -14);
Signal SumNode_Float146Output_667: float (5 downto -14);
Signal ProductNode_Float521Output_668: float (5 downto -14);
Signal ProductNode_Float522weight : float ( 5 downto -14 ) := to_float (0.919167,5,14);

Signal ProductNode_Float522Output_669: float (5 downto -14);
Signal ProductNode_Float523weight : float ( 5 downto -14 ) := to_float (0.781132,5,14);

Signal ProductNode_Float523Output_670: float (5 downto -14);
Signal SumNode_Float147Output_671: float (5 downto -14);
Signal ProductNode_Float524Output_672: float (5 downto -14);
Signal ProductNode_Float525weight : float ( 5 downto -14 ) := to_float (0.970921,5,14);

Signal ProductNode_Float525Output_673: float (5 downto -14);
Signal ProductNode_Float526weight : float ( 5 downto -14 ) := to_float (0.672140,5,14);

Signal ProductNode_Float526Output_674: float (5 downto -14);
Signal SumNode_Float148Output_675: float (5 downto -14);
Signal ProductNode_Float527Output_676: float (5 downto -14);
Signal ProductNode_Float528weight : float ( 5 downto -14 ) := to_float (0.989270,5,14);

Signal ProductNode_Float528Output_677: float (5 downto -14);
Signal ProductNode_Float529weight : float ( 5 downto -14 ) := to_float (0.966381,5,14);

Signal ProductNode_Float529Output_678: float (5 downto -14);
Signal ProductNode_Float530weight : float ( 5 downto -14 ) := to_float (0.690672,5,14);

Signal ProductNode_Float530Output_679: float (5 downto -14);
Signal SumNode_Float149Output_680: float (5 downto -14);
Signal ProductNode_Float531Output_681: float (5 downto -14);
Signal ProductNode_Float532weight : float ( 5 downto -14 ) := to_float (0.853307,5,14);

Signal ProductNode_Float532Output_682: float (5 downto -14);
Signal ProductNode_Float533weight : float ( 5 downto -14 ) := to_float (0.886527,5,14);

Signal ProductNode_Float533Output_683: float (5 downto -14);
Signal SumNode_Float150Output_684: float (5 downto -14);
Signal ProductNode_Float534Output_685: float (5 downto -14);
Signal ProductNode_Float535weight : float ( 5 downto -14 ) := to_float (0.554692,5,14);

Signal ProductNode_Float535Output_686: float (5 downto -14);
Signal ProductNode_Float536weight : float ( 5 downto -14 ) := to_float (0.941870,5,14);

Signal ProductNode_Float536Output_687: float (5 downto -14);
Signal ProductNode_Float537weight : float ( 5 downto -14 ) := to_float (0.763101,5,14);

Signal ProductNode_Float537Output_688: float (5 downto -14);
Signal SumNode_Float151Output_689: float (5 downto -14);
Signal ProductNode_Float538Output_690: float (5 downto -14);
Signal SumNode_Float152Output_691: float (5 downto -14);
Signal ProductNode_Float539Output_692: float (5 downto -14);
Signal ProductNode_Float540weight : float ( 5 downto -14 ) := to_float (0.840616,5,14);

Signal ProductNode_Float540Output_693: float (5 downto -14);
Signal ProductNode_Float541weight : float ( 5 downto -14 ) := to_float (0.817897,5,14);

Signal ProductNode_Float541Output_694: float (5 downto -14);
Signal ProductNode_Float542weight : float ( 5 downto -14 ) := to_float (0.912886,5,14);

Signal ProductNode_Float542Output_695: float (5 downto -14);
Signal SumNode_Float153Output_696: float (5 downto -14);
Signal ProductNode_Float543Output_697: float (5 downto -14);
Signal ProductNode_Float544weight : float ( 5 downto -14 ) := to_float (0.976301,5,14);

Signal ProductNode_Float544Output_698: float (5 downto -14);
Signal ProductNode_Float545weight : float ( 5 downto -14 ) := to_float (0.909585,5,14);

Signal ProductNode_Float545Output_699: float (5 downto -14);
Signal ProductNode_Float546weight : float ( 5 downto -14 ) := to_float (0.822920,5,14);

Signal ProductNode_Float546Output_700: float (5 downto -14);
Signal SumNode_Float154Output_701: float (5 downto -14);
Signal ProductNode_Float547Output_702: float (5 downto -14);
Signal ProductNode_Float548weight : float ( 5 downto -14 ) := to_float (0.731617,5,14);

Signal ProductNode_Float548Output_703: float (5 downto -14);
Signal ProductNode_Float549weight : float ( 5 downto -14 ) := to_float (0.954043,5,14);

Signal ProductNode_Float549Output_704: float (5 downto -14);
Signal SumNode_Float155Output_705: float (5 downto -14);
Signal ProductNode_Float550Output_706: float (5 downto -14);
Signal ProductNode_Float551weight : float ( 5 downto -14 ) := to_float (0.646579,5,14);

Signal ProductNode_Float551Output_707: float (5 downto -14);
Signal ProductNode_Float552weight : float ( 5 downto -14 ) := to_float (0.790147,5,14);

Signal ProductNode_Float552Output_708: float (5 downto -14);
Signal ProductNode_Float553weight : float ( 5 downto -14 ) := to_float (0.929014,5,14);

Signal ProductNode_Float553Output_709: float (5 downto -14);
Signal SumNode_Float156Output_710: float (5 downto -14);
Signal ProductNode_Float554Output_711: float (5 downto -14);
Signal SumNode_Float157Output_712: float (5 downto -14);
Signal ProductNode_Float555Output_713: float (5 downto -14);
Signal ProductNode_Float556weight : float ( 5 downto -14 ) := to_float (0.896858,5,14);

Signal ProductNode_Float556Output_714: float (5 downto -14);
Signal SumNode_Float158Output_715: float (5 downto -14);
Signal ProductNode_Float557Output_716: float (5 downto -14);
Signal ProductNode_Float558weight : float ( 5 downto -14 ) := to_float (0.750079,5,14);

Signal ProductNode_Float558Output_717: float (5 downto -14);
Signal ProductNode_Float559weight : float ( 5 downto -14 ) := to_float (0.947231,5,14);

Signal ProductNode_Float559Output_718: float (5 downto -14);
Signal SumNode_Float159Output_719: float (5 downto -14);
Signal ProductNode_Float560Output_720: float (5 downto -14);
Signal ProductNode_Float561weight : float ( 5 downto -14 ) := to_float (0.807766,5,14);

Signal ProductNode_Float561Output_721: float (5 downto -14);
Signal ProductNode_Float562weight : float ( 5 downto -14 ) := to_float (0.825885,5,14);

Signal ProductNode_Float562Output_722: float (5 downto -14);
Signal ProductNode_Float563weight : float ( 5 downto -14 ) := to_float (0.617466,5,14);

Signal ProductNode_Float563Output_723: float (5 downto -14);
Signal ProductNode_Float564weight : float ( 5 downto -14 ) := to_float (0.981367,5,14);

Signal ProductNode_Float564Output_724: float (5 downto -14);
Signal SumNode_Float160Output_725: float (5 downto -14);
Signal ProductNode_Float565Output_726: float (5 downto -14);
Signal ProductNode_Float566weight : float ( 5 downto -14 ) := to_float (0.919167,5,14);

Signal ProductNode_Float566Output_727: float (5 downto -14);
Signal ProductNode_Float567weight : float ( 5 downto -14 ) := to_float (0.933580,5,14);

Signal ProductNode_Float567Output_728: float (5 downto -14);
Signal SumNode_Float161Output_729: float (5 downto -14);
Signal ProductNode_Float568Output_730: float (5 downto -14);
Signal SumNode_Float162Output_731: float (5 downto -14);
Signal ProductNode_Float569Output_732: float (5 downto -14);
Signal ProductNode_Float570weight : float ( 5 downto -14 ) := to_float (0.776577,5,14);

Signal ProductNode_Float570Output_733: float (5 downto -14);
Signal SumNode_Float163Output_734: float (5 downto -14);
Signal ProductNode_Float571Output_735: float (5 downto -14);
Signal SumNode_Float164Output_736: float (5 downto -14);
Signal ProductNode_Float572Output_737: float (5 downto -14);
Signal ProductNode_Float573weight : float ( 5 downto -14 ) := to_float (0.848299,5,14);

Signal ProductNode_Float573Output_738: float (5 downto -14);
Signal ProductNode_Float574weight : float ( 5 downto -14 ) := to_float (0.895308,5,14);

Signal ProductNode_Float574Output_739: float (5 downto -14);
Signal ProductNode_Float575weight : float ( 5 downto -14 ) := to_float (0.842608,5,14);

Signal ProductNode_Float575Output_740: float (5 downto -14);
Signal SumNode_Float165Output_741: float (5 downto -14);
Signal ProductNode_Float576Output_742: float (5 downto -14);
Signal ProductNode_Float577weight : float ( 5 downto -14 ) := to_float (0.870697,5,14);

Signal ProductNode_Float577Output_743: float (5 downto -14);
Signal ProductNode_Float578weight : float ( 5 downto -14 ) := to_float (0.945793,5,14);

Signal ProductNode_Float578Output_744: float (5 downto -14);
Signal ProductNode_Float579weight : float ( 5 downto -14 ) := to_float (0.954870,5,14);

Signal ProductNode_Float579Output_745: float (5 downto -14);
Signal ProductNode_Float580weight : float ( 5 downto -14 ) := to_float (0.870404,5,14);

Signal ProductNode_Float580Output_746: float (5 downto -14);
Signal ProductNode_Float581weight : float ( 5 downto -14 ) := to_float (0.780732,5,14);

Signal ProductNode_Float581Output_747: float (5 downto -14);
Signal ProductNode_Float582weight : float ( 5 downto -14 ) := to_float (0.810846,5,14);

Signal ProductNode_Float582Output_748: float (5 downto -14);
Signal SumNode_Float166Output_749: float (5 downto -14);
Signal ProductNode_Float583Output_750: float (5 downto -14);
Signal ProductNode_Float584weight : float ( 5 downto -14 ) := to_float (0.531606,5,14);

Signal ProductNode_Float584Output_751: float (5 downto -14);
Signal ProductNode_Float585weight : float ( 5 downto -14 ) := to_float (0.669241,5,14);

Signal ProductNode_Float585Output_752: float (5 downto -14);
Signal ProductNode_Float586weight : float ( 5 downto -14 ) := to_float (0.971580,5,14);

Signal ProductNode_Float586Output_753: float (5 downto -14);
Signal SumNode_Float167Output_754: float (5 downto -14);
Signal ProductNode_Float587Output_755: float (5 downto -14);
Signal ProductNode_Float588weight : float ( 5 downto -14 ) := to_float (0.870697,5,14);

Signal ProductNode_Float588Output_756: float (5 downto -14);
Signal ProductNode_Float589weight : float ( 5 downto -14 ) := to_float (0.753690,5,14);

Signal ProductNode_Float589Output_757: float (5 downto -14);
Signal ProductNode_Float590weight : float ( 5 downto -14 ) := to_float (0.774480,5,14);

Signal ProductNode_Float590Output_758: float (5 downto -14);
Signal ProductNode_Float591weight : float ( 5 downto -14 ) := to_float (0.870404,5,14);

Signal ProductNode_Float591Output_759: float (5 downto -14);
Signal ProductNode_Float592weight : float ( 5 downto -14 ) := to_float (0.933776,5,14);

Signal ProductNode_Float592Output_760: float (5 downto -14);
Signal ProductNode_Float593weight : float ( 5 downto -14 ) := to_float (0.660973,5,14);

Signal ProductNode_Float593Output_761: float (5 downto -14);
Signal SumNode_Float168Output_762: float (5 downto -14);
Signal ProductNode_Float594Output_763: float (5 downto -14);
Signal ProductNode_Float595weight : float ( 5 downto -14 ) := to_float (0.870862,5,14);

Signal ProductNode_Float595Output_764: float (5 downto -14);
Signal SumNode_Float169Output_765: float (5 downto -14);
Signal ProductNode_Float596Output_766: float (5 downto -14);
Signal ProductNode_Float597weight : float ( 5 downto -14 ) := to_float (0.850730,5,14);

Signal ProductNode_Float597Output_767: float (5 downto -14);
Signal ProductNode_Float598weight : float ( 5 downto -14 ) := to_float (0.890735,5,14);

Signal ProductNode_Float598Output_768: float (5 downto -14);
Signal ProductNode_Float599weight : float ( 5 downto -14 ) := to_float (0.689002,5,14);

Signal ProductNode_Float599Output_769: float (5 downto -14);
Signal ProductNode_Float600weight : float ( 5 downto -14 ) := to_float (0.966814,5,14);

Signal ProductNode_Float600Output_770: float (5 downto -14);
Signal SumNode_Float170Output_771: float (5 downto -14);
Signal ProductNode_Float601Output_772: float (5 downto -14);
Signal ProductNode_Float602weight : float ( 5 downto -14 ) := to_float (0.551341,5,14);

Signal ProductNode_Float602Output_773: float (5 downto -14);
Signal ProductNode_Float603weight : float ( 5 downto -14 ) := to_float (0.795357,5,14);

Signal ProductNode_Float603Output_774: float (5 downto -14);
Signal ProductNode_Float604weight : float ( 5 downto -14 ) := to_float (0.746308,5,14);

Signal ProductNode_Float604Output_775: float (5 downto -14);
Signal ProductNode_Float605weight : float ( 5 downto -14 ) := to_float (0.989597,5,14);

Signal ProductNode_Float605Output_776: float (5 downto -14);
Signal ProductNode_Float606weight : float ( 5 downto -14 ) := to_float (0.577708,5,14);

Signal ProductNode_Float606Output_777: float (5 downto -14);
Signal ProductNode_Float607weight : float ( 5 downto -14 ) := to_float (0.618274,5,14);

Signal ProductNode_Float607Output_778: float (5 downto -14);
Signal SumNode_Float171Output_779: float (5 downto -14);
Signal ProductNode_Float608Output_780: float (5 downto -14);
Signal ProductNode_Float609weight : float ( 5 downto -14 ) := to_float (0.735141,5,14);

Signal ProductNode_Float609Output_781: float (5 downto -14);
Signal ProductNode_Float610weight : float ( 5 downto -14 ) := to_float (0.495915,5,14);

Signal ProductNode_Float610Output_782: float (5 downto -14);
Signal ProductNode_Float611weight : float ( 5 downto -14 ) := to_float (0.993928,5,14);

Signal ProductNode_Float611Output_783: float (5 downto -14);
Signal SumNode_Float172Output_784: float (5 downto -14);
Signal ProductNode_Float612Output_785: float (5 downto -14);
Signal ProductNode_Float613weight : float ( 5 downto -14 ) := to_float (0.551341,5,14);

Signal ProductNode_Float613Output_786: float (5 downto -14);
Signal ProductNode_Float614weight : float ( 5 downto -14 ) := to_float (0.926235,5,14);

Signal ProductNode_Float614Output_787: float (5 downto -14);
Signal ProductNode_Float615weight : float ( 5 downto -14 ) := to_float (0.616494,5,14);

Signal ProductNode_Float615Output_788: float (5 downto -14);
Signal ProductNode_Float616weight : float ( 5 downto -14 ) := to_float (0.989597,5,14);

Signal ProductNode_Float616Output_789: float (5 downto -14);
Signal ProductNode_Float617weight : float ( 5 downto -14 ) := to_float (0.986786,5,14);

Signal ProductNode_Float617Output_790: float (5 downto -14);
Signal ProductNode_Float618weight : float ( 5 downto -14 ) := to_float (0.464416,5,14);

Signal ProductNode_Float618Output_791: float (5 downto -14);
Signal SumNode_Float173Output_792: float (5 downto -14);
Signal ProductNode_Float619Output_793: float (5 downto -14);
Signal ProductNode_Float620weight : float ( 5 downto -14 ) := to_float (0.938375,5,14);

Signal ProductNode_Float620Output_794: float (5 downto -14);
Signal SumNode_Float174Output_795: float (5 downto -14);
Signal ProductNode_Float621Output_796: float (5 downto -14);
Signal ProductNode_Float622weight : float ( 5 downto -14 ) := to_float (0.635106,5,14);

Signal ProductNode_Float622Output_797: float (5 downto -14);
Signal SumNode_Float175Output_798: float (5 downto -14);
Signal ProductNode_Float623Output_799: float (5 downto -14);
Signal ProductNode_Float624weight : float ( 5 downto -14 ) := to_float (0.969587,5,14);

Signal ProductNode_Float624Output_800: float (5 downto -14);
Signal ProductNode_Float625weight : float ( 5 downto -14 ) := to_float (0.848299,5,14);

Signal ProductNode_Float625Output_801: float (5 downto -14);
Signal ProductNode_Float626weight : float ( 5 downto -14 ) := to_float (0.562709,5,14);

Signal ProductNode_Float626Output_802: float (5 downto -14);
Signal ProductNode_Float627weight : float ( 5 downto -14 ) := to_float (0.988453,5,14);

Signal ProductNode_Float627Output_803: float (5 downto -14);
Signal SumNode_Float176Output_804: float (5 downto -14);
Signal ProductNode_Float628Output_805: float (5 downto -14);
Signal ProductNode_Float629weight : float ( 5 downto -14 ) := to_float (0.870697,5,14);

Signal ProductNode_Float629Output_806: float (5 downto -14);
Signal ProductNode_Float630weight : float ( 5 downto -14 ) := to_float (0.945793,5,14);

Signal ProductNode_Float630Output_807: float (5 downto -14);
Signal ProductNode_Float631weight : float ( 5 downto -14 ) := to_float (0.729204,5,14);

Signal ProductNode_Float631Output_808: float (5 downto -14);
Signal ProductNode_Float632weight : float ( 5 downto -14 ) := to_float (0.870404,5,14);

Signal ProductNode_Float632Output_809: float (5 downto -14);
Signal ProductNode_Float633weight : float ( 5 downto -14 ) := to_float (0.780732,5,14);

Signal ProductNode_Float633Output_810: float (5 downto -14);
Signal ProductNode_Float634weight : float ( 5 downto -14 ) := to_float (0.917308,5,14);

Signal ProductNode_Float634Output_811: float (5 downto -14);
Signal SumNode_Float177Output_812: float (5 downto -14);
Signal ProductNode_Float635Output_813: float (5 downto -14);
Signal ProductNode_Float636weight : float ( 5 downto -14 ) := to_float (0.631626,5,14);

Signal ProductNode_Float636Output_814: float (5 downto -14);
Signal ProductNode_Float637weight : float ( 5 downto -14 ) := to_float (0.453222,5,14);

Signal ProductNode_Float637Output_815: float (5 downto -14);
Signal ProductNode_Float638weight : float ( 5 downto -14 ) := to_float (0.996146,5,14);

Signal ProductNode_Float638Output_816: float (5 downto -14);
Signal SumNode_Float178Output_817: float (5 downto -14);
Signal ProductNode_Float639Output_818: float (5 downto -14);
Signal ProductNode_Float640weight : float ( 5 downto -14 ) := to_float (0.870697,5,14);

Signal ProductNode_Float640Output_819: float (5 downto -14);
Signal ProductNode_Float641weight : float ( 5 downto -14 ) := to_float (0.753690,5,14);

Signal ProductNode_Float641Output_820: float (5 downto -14);
Signal ProductNode_Float642weight : float ( 5 downto -14 ) := to_float (0.936763,5,14);

Signal ProductNode_Float642Output_821: float (5 downto -14);
Signal ProductNode_Float643weight : float ( 5 downto -14 ) := to_float (0.870404,5,14);

Signal ProductNode_Float643Output_822: float (5 downto -14);
Signal ProductNode_Float644weight : float ( 5 downto -14 ) := to_float (0.933776,5,14);

Signal ProductNode_Float644Output_823: float (5 downto -14);
Signal ProductNode_Float645weight : float ( 5 downto -14 ) := to_float (0.973389,5,14);

Signal ProductNode_Float645Output_824: float (5 downto -14);
Signal SumNode_Float179Output_825: float (5 downto -14);
Signal ProductNode_Float646Output_826: float (5 downto -14);
Signal ProductNode_Float647weight : float ( 5 downto -14 ) := to_float (0.912549,5,14);

Signal ProductNode_Float647Output_827: float (5 downto -14);
Signal SumNode_Float180Output_828: float (5 downto -14);
Signal ProductNode_Float648Output_829: float (5 downto -14);
Signal ProductNode_Float649weight : float ( 5 downto -14 ) := to_float (0.658116,5,14);

Signal ProductNode_Float649Output_830: float (5 downto -14);
Signal ProductNode_Float650weight : float ( 5 downto -14 ) := to_float (0.890735,5,14);

Signal ProductNode_Float650Output_831: float (5 downto -14);
Signal ProductNode_Float651weight : float ( 5 downto -14 ) := to_float (0.382644,5,14);

Signal ProductNode_Float651Output_832: float (5 downto -14);
Signal ProductNode_Float652weight : float ( 5 downto -14 ) := to_float (0.998354,5,14);

Signal ProductNode_Float652Output_833: float (5 downto -14);
Signal SumNode_Float181Output_834: float (5 downto -14);
Signal ProductNode_Float653Output_835: float (5 downto -14);
Signal ProductNode_Float654weight : float ( 5 downto -14 ) := to_float (0.551341,5,14);

Signal ProductNode_Float654Output_836: float (5 downto -14);
Signal ProductNode_Float655weight : float ( 5 downto -14 ) := to_float (0.795357,5,14);

Signal ProductNode_Float655Output_837: float (5 downto -14);
Signal ProductNode_Float656weight : float ( 5 downto -14 ) := to_float (0.948695,5,14);

Signal ProductNode_Float656Output_838: float (5 downto -14);
Signal ProductNode_Float657weight : float ( 5 downto -14 ) := to_float (0.989597,5,14);

Signal ProductNode_Float657Output_839: float (5 downto -14);
Signal ProductNode_Float658weight : float ( 5 downto -14 ) := to_float (0.577708,5,14);

Signal ProductNode_Float658Output_840: float (5 downto -14);
Signal ProductNode_Float659weight : float ( 5 downto -14 ) := to_float (0.981240,5,14);

Signal ProductNode_Float659Output_841: float (5 downto -14);
Signal SumNode_Float182Output_842: float (5 downto -14);
Signal ProductNode_Float660Output_843: float (5 downto -14);
Signal ProductNode_Float661weight : float ( 5 downto -14 ) := to_float (0.712179,5,14);

Signal ProductNode_Float661Output_844: float (5 downto -14);
Signal ProductNode_Float662weight : float ( 5 downto -14 ) := to_float (0.336149,5,14);

Signal ProductNode_Float662Output_845: float (5 downto -14);
Signal ProductNode_Float663weight : float ( 5 downto -14 ) := to_float (0.999140,5,14);

Signal ProductNode_Float663Output_846: float (5 downto -14);
Signal SumNode_Float183Output_847: float (5 downto -14);
Signal ProductNode_Float664Output_848: float (5 downto -14);
Signal ProductNode_Float665weight : float ( 5 downto -14 ) := to_float (0.551341,5,14);

Signal ProductNode_Float665Output_849: float (5 downto -14);
Signal ProductNode_Float666weight : float ( 5 downto -14 ) := to_float (0.926235,5,14);

Signal ProductNode_Float666Output_850: float (5 downto -14);
Signal ProductNode_Float667weight : float ( 5 downto -14 ) := to_float (0.981519,5,14);

Signal ProductNode_Float667Output_851: float (5 downto -14);
Signal ProductNode_Float668weight : float ( 5 downto -14 ) := to_float (0.989597,5,14);

Signal ProductNode_Float668Output_852: float (5 downto -14);
Signal ProductNode_Float669weight : float ( 5 downto -14 ) := to_float (0.986786,5,14);

Signal ProductNode_Float669Output_853: float (5 downto -14);
Signal ProductNode_Float670weight : float ( 5 downto -14 ) := to_float (0.995641,5,14);

Signal ProductNode_Float670Output_854: float (5 downto -14);
Signal SumNode_Float184Output_855: float (5 downto -14);
Signal ProductNode_Float671Output_856: float (5 downto -14);
Signal ProductNode_Float672weight : float ( 5 downto -14 ) := to_float (0.972670,5,14);

Signal ProductNode_Float672Output_857: float (5 downto -14);
Signal SumNode_Float185Output_858: float (5 downto -14);
Signal ProductNode_Float673Output_859: float (5 downto -14);
Signal ProductNode_Float674weight : float ( 5 downto -14 ) := to_float (0.531350,5,14);

Signal ProductNode_Float674Output_860: float (5 downto -14);
Signal SumNode_Float186Output_861: float (5 downto -14);
Signal ProductNode_Float675Output_862: float (5 downto -14);
Signal ProductNode_Float676weight : float ( 5 downto -14 ) := to_float (0.913608,5,14);

Signal ProductNode_Float676Output_863: float (5 downto -14);
Signal SumNode_Float187Output_864: float (5 downto -14);
Signal ProductNode_Float677Output_865: float (5 downto -14);
Signal ProductNode_Float678weight : float ( 5 downto -14 ) := to_float (0.965849,5,14);

Signal ProductNode_Float678Output_866: float (5 downto -14);
Signal ProductNode_Float679weight : float ( 5 downto -14 ) := to_float (0.692695,5,14);

Signal ProductNode_Float679Output_867: float (5 downto -14);
Signal SumNode_Float188Output_868: float (5 downto -14);
Signal ProductNode_Float680Output_869: float (5 downto -14);
Signal ProductNode_Float681weight : float ( 5 downto -14 ) := to_float (0.880399,5,14);

Signal ProductNode_Float681Output_870: float (5 downto -14);
Signal ProductNode_Float682weight : float ( 5 downto -14 ) := to_float (0.997554,5,14);

Signal ProductNode_Float682Output_871: float (5 downto -14);
Signal ProductNode_Float683weight : float ( 5 downto -14 ) := to_float (0.414069,5,14);

Signal ProductNode_Float683Output_872: float (5 downto -14);
Signal SumNode_Float189Output_873: float (5 downto -14);
Signal ProductNode_Float684Output_874: float (5 downto -14);
Signal ProductNode_Float685weight : float ( 5 downto -14 ) := to_float (0.919660,5,14);

Signal ProductNode_Float685Output_875: float (5 downto -14);
Signal ProductNode_Float686weight : float ( 5 downto -14 ) := to_float (0.806938,5,14);

Signal ProductNode_Float686Output_876: float (5 downto -14);
Signal SumNode_Float190Output_877: float (5 downto -14);
Signal ProductNode_Float687Output_878: float (5 downto -14);
Signal ProductNode_Float688weight : float ( 5 downto -14 ) := to_float (0.860235,5,14);

Signal ProductNode_Float688Output_879: float (5 downto -14);
Signal ProductNode_Float689weight : float ( 5 downto -14 ) := to_float (0.989739,5,14);

Signal ProductNode_Float689Output_880: float (5 downto -14);
Signal ProductNode_Float690weight : float ( 5 downto -14 ) := to_float (0.549861,5,14);

Signal ProductNode_Float690Output_881: float (5 downto -14);
Signal SumNode_Float191Output_882: float (5 downto -14);
Signal ProductNode_Float691Output_883: float (5 downto -14);
Signal SumNode_Float192Output_884: float (5 downto -14);
Signal ProductNode_Float692Output_885: float (5 downto -14);
Signal ProductNode_Float693weight : float ( 5 downto -14 ) := to_float (0.984104,5,14);

Signal ProductNode_Float693Output_886: float (5 downto -14);
Signal ProductNode_Float694weight : float ( 5 downto -14 ) := to_float (0.793165,5,14);

Signal ProductNode_Float694Output_887: float (5 downto -14);
Signal ProductNode_Float695weight : float ( 5 downto -14 ) := to_float (0.927417,5,14);

Signal ProductNode_Float695Output_888: float (5 downto -14);
Signal SumNode_Float193Output_889: float (5 downto -14);
Signal ProductNode_Float696Output_890: float (5 downto -14);
Signal ProductNode_Float697weight : float ( 5 downto -14 ) := to_float (0.726095,5,14);

Signal ProductNode_Float697Output_891: float (5 downto -14);
Signal ProductNode_Float698weight : float ( 5 downto -14 ) := to_float (0.988880,5,14);

Signal ProductNode_Float698Output_892: float (5 downto -14);
Signal ProductNode_Float699weight : float ( 5 downto -14 ) := to_float (0.558577,5,14);

Signal ProductNode_Float699Output_893: float (5 downto -14);
Signal SumNode_Float194Output_894: float (5 downto -14);
Signal ProductNode_Float700Output_895: float (5 downto -14);
Signal ProductNode_Float701weight : float ( 5 downto -14 ) := to_float (0.649155,5,14);

Signal ProductNode_Float701Output_896: float (5 downto -14);
Signal ProductNode_Float702weight : float ( 5 downto -14 ) := to_float (0.975801,5,14);

Signal ProductNode_Float702Output_897: float (5 downto -14);
Signal SumNode_Float195Output_898: float (5 downto -14);
Signal ProductNode_Float703Output_899: float (5 downto -14);
Signal ProductNode_Float704weight : float ( 5 downto -14 ) := to_float (0.955917,5,14);

Signal ProductNode_Float704Output_900: float (5 downto -14);
Signal ProductNode_Float705weight : float ( 5 downto -14 ) := to_float (0.985013,5,14);

Signal ProductNode_Float705Output_901: float (5 downto -14);
Signal ProductNode_Float706weight : float ( 5 downto -14 ) := to_float (0.592017,5,14);

Signal ProductNode_Float706Output_902: float (5 downto -14);
Signal SumNode_Float196Output_903: float (5 downto -14);
Signal ProductNode_Float707Output_904: float (5 downto -14);
Signal SumNode_Float197Output_905: float (5 downto -14);
Signal ProductNode_Float708Output_906: float (5 downto -14);
Signal ProductNode_Float709weight : float ( 5 downto -14 ) := to_float (0.598812,5,14);

Signal ProductNode_Float709Output_907: float (5 downto -14);
Signal SumNode_Float198Output_908: float (5 downto -14);
Signal ProductNode_Float710Output_909: float (5 downto -14);
Signal ProductNode_Float711weight : float ( 5 downto -14 ) := to_float (0.927615,5,14);

Signal ProductNode_Float711Output_910: float (5 downto -14);
Signal ProductNode_Float712weight : float ( 5 downto -14 ) := to_float (0.792795,5,14);

Signal ProductNode_Float712Output_911: float (5 downto -14);
Signal SumNode_Float199Output_912: float (5 downto -14);
Signal ProductNode_Float713Output_913: float (5 downto -14);
Signal ProductNode_Float714weight : float ( 5 downto -14 ) := to_float (0.907425,5,14);

Signal ProductNode_Float714Output_914: float (5 downto -14);
Signal ProductNode_Float715weight : float ( 5 downto -14 ) := to_float (0.948402,5,14);

Signal ProductNode_Float715Output_915: float (5 downto -14);
Signal ProductNode_Float716weight : float ( 5 downto -14 ) := to_float (0.838940,5,14);

Signal ProductNode_Float716Output_916: float (5 downto -14);
Signal ProductNode_Float717weight : float ( 5 downto -14 ) := to_float (0.898142,5,14);

Signal ProductNode_Float717Output_917: float (5 downto -14);
Signal SumNode_Float200Output_918: float (5 downto -14);
Signal ProductNode_Float718Output_919: float (5 downto -14);
Signal ProductNode_Float719weight : float ( 5 downto -14 ) := to_float (0.826105,5,14);

Signal ProductNode_Float719Output_920: float (5 downto -14);
Signal ProductNode_Float720weight : float ( 5 downto -14 ) := to_float (0.838083,5,14);

Signal ProductNode_Float720Output_921: float (5 downto -14);
Signal SumNode_Float201Output_922: float (5 downto -14);
Signal ProductNode_Float721Output_923: float (5 downto -14);
Signal ProductNode_Float722weight : float ( 5 downto -14 ) := to_float (0.965849,5,14);

Signal ProductNode_Float722Output_924: float (5 downto -14);
Signal ProductNode_Float723weight : float ( 5 downto -14 ) := to_float (0.692695,5,14);

Signal ProductNode_Float723Output_925: float (5 downto -14);
Signal SumNode_Float202Output_926: float (5 downto -14);
Signal ProductNode_Float724Output_927: float (5 downto -14);
Signal ProductNode_Float725weight : float ( 5 downto -14 ) := to_float (0.880399,5,14);

Signal ProductNode_Float725Output_928: float (5 downto -14);
Signal ProductNode_Float726weight : float ( 5 downto -14 ) := to_float (0.997554,5,14);

Signal ProductNode_Float726Output_929: float (5 downto -14);
Signal ProductNode_Float727weight : float ( 5 downto -14 ) := to_float (0.414069,5,14);

Signal ProductNode_Float727Output_930: float (5 downto -14);
Signal SumNode_Float203Output_931: float (5 downto -14);
Signal ProductNode_Float728Output_932: float (5 downto -14);
Signal ProductNode_Float729weight : float ( 5 downto -14 ) := to_float (0.919660,5,14);

Signal ProductNode_Float729Output_933: float (5 downto -14);
Signal ProductNode_Float730weight : float ( 5 downto -14 ) := to_float (0.806938,5,14);

Signal ProductNode_Float730Output_934: float (5 downto -14);
Signal SumNode_Float204Output_935: float (5 downto -14);
Signal ProductNode_Float731Output_936: float (5 downto -14);
Signal ProductNode_Float732weight : float ( 5 downto -14 ) := to_float (0.860235,5,14);

Signal ProductNode_Float732Output_937: float (5 downto -14);
Signal ProductNode_Float733weight : float ( 5 downto -14 ) := to_float (0.989739,5,14);

Signal ProductNode_Float733Output_938: float (5 downto -14);
Signal ProductNode_Float734weight : float ( 5 downto -14 ) := to_float (0.549861,5,14);

Signal ProductNode_Float734Output_939: float (5 downto -14);
Signal SumNode_Float205Output_940: float (5 downto -14);
Signal ProductNode_Float735Output_941: float (5 downto -14);
Signal SumNode_Float206Output_942: float (5 downto -14);
Signal ProductNode_Float736Output_943: float (5 downto -14);
Signal ProductNode_Float737weight : float ( 5 downto -14 ) := to_float (0.932937,5,14);

Signal ProductNode_Float737Output_944: float (5 downto -14);
Signal ProductNode_Float738weight : float ( 5 downto -14 ) := to_float (0.793165,5,14);

Signal ProductNode_Float738Output_945: float (5 downto -14);
Signal ProductNode_Float739weight : float ( 5 downto -14 ) := to_float (0.927417,5,14);

Signal ProductNode_Float739Output_946: float (5 downto -14);
Signal SumNode_Float207Output_947: float (5 downto -14);
Signal ProductNode_Float740Output_948: float (5 downto -14);
Signal ProductNode_Float741weight : float ( 5 downto -14 ) := to_float (0.726095,5,14);

Signal ProductNode_Float741Output_949: float (5 downto -14);
Signal ProductNode_Float742weight : float ( 5 downto -14 ) := to_float (0.988880,5,14);

Signal ProductNode_Float742Output_950: float (5 downto -14);
Signal ProductNode_Float743weight : float ( 5 downto -14 ) := to_float (0.558577,5,14);

Signal ProductNode_Float743Output_951: float (5 downto -14);
Signal SumNode_Float208Output_952: float (5 downto -14);
Signal ProductNode_Float744Output_953: float (5 downto -14);
Signal ProductNode_Float745weight : float ( 5 downto -14 ) := to_float (0.649155,5,14);

Signal ProductNode_Float745Output_954: float (5 downto -14);
Signal ProductNode_Float746weight : float ( 5 downto -14 ) := to_float (0.975801,5,14);

Signal ProductNode_Float746Output_955: float (5 downto -14);
Signal SumNode_Float209Output_956: float (5 downto -14);
Signal ProductNode_Float747Output_957: float (5 downto -14);
Signal ProductNode_Float748weight : float ( 5 downto -14 ) := to_float (0.955917,5,14);

Signal ProductNode_Float748Output_958: float (5 downto -14);
Signal ProductNode_Float749weight : float ( 5 downto -14 ) := to_float (0.985013,5,14);

Signal ProductNode_Float749Output_959: float (5 downto -14);
Signal ProductNode_Float750weight : float ( 5 downto -14 ) := to_float (0.592017,5,14);

Signal ProductNode_Float750Output_960: float (5 downto -14);
Signal SumNode_Float210Output_961: float (5 downto -14);
Signal ProductNode_Float751Output_962: float (5 downto -14);
Signal SumNode_Float211Output_963: float (5 downto -14);
Signal ProductNode_Float752Output_964: float (5 downto -14);
Signal ProductNode_Float753weight : float ( 5 downto -14 ) := to_float (0.782438,5,14);

Signal ProductNode_Float753Output_965: float (5 downto -14);
Signal SumNode_Float212Output_966: float (5 downto -14);
Signal ProductNode_Float754Output_967: float (5 downto -14);
Signal ProductNode_Float755weight : float ( 5 downto -14 ) := to_float (0.750079,5,14);

Signal ProductNode_Float755Output_968: float (5 downto -14);
Signal ProductNode_Float756weight : float ( 5 downto -14 ) := to_float (0.947231,5,14);

Signal ProductNode_Float756Output_969: float (5 downto -14);
Signal SumNode_Float213Output_970: float (5 downto -14);
Signal ProductNode_Float757Output_971: float (5 downto -14);
Signal ProductNode_Float758weight : float ( 5 downto -14 ) := to_float (0.907425,5,14);

Signal ProductNode_Float758Output_972: float (5 downto -14);
Signal ProductNode_Float759weight : float ( 5 downto -14 ) := to_float (0.747070,5,14);

Signal ProductNode_Float759Output_973: float (5 downto -14);
Signal ProductNode_Float760weight : float ( 5 downto -14 ) := to_float (0.617466,5,14);

Signal ProductNode_Float760Output_974: float (5 downto -14);
Signal ProductNode_Float761weight : float ( 5 downto -14 ) := to_float (0.981367,5,14);

Signal ProductNode_Float761Output_975: float (5 downto -14);
Signal SumNode_Float214Output_976: float (5 downto -14);
Signal ProductNode_Float762Output_977: float (5 downto -14);
Signal ProductNode_Float763weight : float ( 5 downto -14 ) := to_float (0.826105,5,14);

Signal ProductNode_Float763Output_978: float (5 downto -14);
Signal ProductNode_Float764weight : float ( 5 downto -14 ) := to_float (0.898792,5,14);

Signal ProductNode_Float764Output_979: float (5 downto -14);
Signal SumNode_Float215Output_980: float (5 downto -14);
Signal ProductNode_Float765Output_981: float (5 downto -14);
Signal SumNode_Float216Output_982: float (5 downto -14);
Signal ProductNode_Float766Output_983: float (5 downto -14);
Signal ProductNode_Float767weight : float ( 5 downto -14 ) := to_float (0.987852,5,14);

Signal ProductNode_Float767Output_984: float (5 downto -14);
Signal ProductNode_Float768weight : float ( 5 downto -14 ) := to_float (0.965849,5,14);

Signal ProductNode_Float768Output_985: float (5 downto -14);
Signal ProductNode_Float769weight : float ( 5 downto -14 ) := to_float (0.692695,5,14);

Signal ProductNode_Float769Output_986: float (5 downto -14);
Signal SumNode_Float217Output_987: float (5 downto -14);
Signal ProductNode_Float770Output_988: float (5 downto -14);
Signal ProductNode_Float771weight : float ( 5 downto -14 ) := to_float (0.880399,5,14);

Signal ProductNode_Float771Output_989: float (5 downto -14);
Signal ProductNode_Float772weight : float ( 5 downto -14 ) := to_float (0.966381,5,14);

Signal ProductNode_Float772Output_990: float (5 downto -14);
Signal ProductNode_Float773weight : float ( 5 downto -14 ) := to_float (0.690672,5,14);

Signal ProductNode_Float773Output_991: float (5 downto -14);
Signal SumNode_Float218Output_992: float (5 downto -14);
Signal ProductNode_Float774Output_993: float (5 downto -14);
Signal ProductNode_Float775weight : float ( 5 downto -14 ) := to_float (0.919660,5,14);

Signal ProductNode_Float775Output_994: float (5 downto -14);
Signal ProductNode_Float776weight : float ( 5 downto -14 ) := to_float (0.806938,5,14);

Signal ProductNode_Float776Output_995: float (5 downto -14);
Signal SumNode_Float219Output_996: float (5 downto -14);
Signal ProductNode_Float777Output_997: float (5 downto -14);
Signal ProductNode_Float778weight : float ( 5 downto -14 ) := to_float (0.860235,5,14);

Signal ProductNode_Float778Output_998: float (5 downto -14);
Signal ProductNode_Float779weight : float ( 5 downto -14 ) := to_float (0.941870,5,14);

Signal ProductNode_Float779Output_999: float (5 downto -14);
Signal ProductNode_Float780weight : float ( 5 downto -14 ) := to_float (0.763101,5,14);

Signal ProductNode_Float780Output_1000: float (5 downto -14);
Signal SumNode_Float220Output_1001: float (5 downto -14);
Signal ProductNode_Float781Output_1002: float (5 downto -14);
Signal SumNode_Float221Output_1003: float (5 downto -14);
Signal ProductNode_Float782Output_1004: float (5 downto -14);
Signal ProductNode_Float783weight : float ( 5 downto -14 ) := to_float (0.924413,5,14);

Signal ProductNode_Float783Output_1005: float (5 downto -14);
Signal ProductNode_Float784weight : float ( 5 downto -14 ) := to_float (0.793165,5,14);

Signal ProductNode_Float784Output_1006: float (5 downto -14);
Signal ProductNode_Float785weight : float ( 5 downto -14 ) := to_float (0.927417,5,14);

Signal ProductNode_Float785Output_1007: float (5 downto -14);
Signal SumNode_Float222Output_1008: float (5 downto -14);
Signal ProductNode_Float786Output_1009: float (5 downto -14);
Signal ProductNode_Float787weight : float ( 5 downto -14 ) := to_float (0.726095,5,14);

Signal ProductNode_Float787Output_1010: float (5 downto -14);
Signal ProductNode_Float788weight : float ( 5 downto -14 ) := to_float (0.909585,5,14);

Signal ProductNode_Float788Output_1011: float (5 downto -14);
Signal ProductNode_Float789weight : float ( 5 downto -14 ) := to_float (0.822920,5,14);

Signal ProductNode_Float789Output_1012: float (5 downto -14);
Signal SumNode_Float223Output_1013: float (5 downto -14);
Signal ProductNode_Float790Output_1014: float (5 downto -14);
Signal ProductNode_Float791weight : float ( 5 downto -14 ) := to_float (0.649155,5,14);

Signal ProductNode_Float791Output_1015: float (5 downto -14);
Signal ProductNode_Float792weight : float ( 5 downto -14 ) := to_float (0.975801,5,14);

Signal ProductNode_Float792Output_1016: float (5 downto -14);
Signal SumNode_Float224Output_1017: float (5 downto -14);
Signal ProductNode_Float793Output_1018: float (5 downto -14);
Signal ProductNode_Float794weight : float ( 5 downto -14 ) := to_float (0.955917,5,14);

Signal ProductNode_Float794Output_1019: float (5 downto -14);
Signal ProductNode_Float795weight : float ( 5 downto -14 ) := to_float (0.790147,5,14);

Signal ProductNode_Float795Output_1020: float (5 downto -14);
Signal ProductNode_Float796weight : float ( 5 downto -14 ) := to_float (0.929014,5,14);

Signal ProductNode_Float796Output_1021: float (5 downto -14);
Signal SumNode_Float225Output_1022: float (5 downto -14);
Signal ProductNode_Float797Output_1023: float (5 downto -14);
Signal SumNode_Float226Output_1024: float (5 downto -14);
Signal ProductNode_Float798Output_1025: float (5 downto -14);
Signal ProductNode_Float799weight : float ( 5 downto -14 ) := to_float (0.798666,5,14);

Signal ProductNode_Float799Output_1026: float (5 downto -14);
Signal SumNode_Float227Output_1027: float (5 downto -14);
Signal ProductNode_Float800Output_1028: float (5 downto -14);
Signal ProductNode_Float801weight : float ( 5 downto -14 ) := to_float (0.927615,5,14);

Signal ProductNode_Float801Output_1029: float (5 downto -14);
Signal ProductNode_Float802weight : float ( 5 downto -14 ) := to_float (0.792795,5,14);

Signal ProductNode_Float802Output_1030: float (5 downto -14);
Signal SumNode_Float228Output_1031: float (5 downto -14);
Signal ProductNode_Float803Output_1032: float (5 downto -14);
Signal ProductNode_Float804weight : float ( 5 downto -14 ) := to_float (0.807766,5,14);

Signal ProductNode_Float804Output_1033: float (5 downto -14);
Signal ProductNode_Float805weight : float ( 5 downto -14 ) := to_float (0.907576,5,14);

Signal ProductNode_Float805Output_1034: float (5 downto -14);
Signal ProductNode_Float806weight : float ( 5 downto -14 ) := to_float (0.838940,5,14);

Signal ProductNode_Float806Output_1035: float (5 downto -14);
Signal ProductNode_Float807weight : float ( 5 downto -14 ) := to_float (0.898142,5,14);

Signal ProductNode_Float807Output_1036: float (5 downto -14);
Signal SumNode_Float229Output_1037: float (5 downto -14);
Signal ProductNode_Float808Output_1038: float (5 downto -14);
Signal ProductNode_Float809weight : float ( 5 downto -14 ) := to_float (0.919167,5,14);

Signal ProductNode_Float809Output_1039: float (5 downto -14);
Signal ProductNode_Float810weight : float ( 5 downto -14 ) := to_float (0.781132,5,14);

Signal ProductNode_Float810Output_1040: float (5 downto -14);
Signal SumNode_Float230Output_1041: float (5 downto -14);
Signal ProductNode_Float811Output_1042: float (5 downto -14);
Signal ProductNode_Float812weight : float ( 5 downto -14 ) := to_float (0.965849,5,14);

Signal ProductNode_Float812Output_1043: float (5 downto -14);
Signal ProductNode_Float813weight : float ( 5 downto -14 ) := to_float (0.692695,5,14);

Signal ProductNode_Float813Output_1044: float (5 downto -14);
Signal SumNode_Float231Output_1045: float (5 downto -14);
Signal ProductNode_Float814Output_1046: float (5 downto -14);
Signal ProductNode_Float815weight : float ( 5 downto -14 ) := to_float (0.880399,5,14);

Signal ProductNode_Float815Output_1047: float (5 downto -14);
Signal ProductNode_Float816weight : float ( 5 downto -14 ) := to_float (0.966381,5,14);

Signal ProductNode_Float816Output_1048: float (5 downto -14);
Signal ProductNode_Float817weight : float ( 5 downto -14 ) := to_float (0.690672,5,14);

Signal ProductNode_Float817Output_1049: float (5 downto -14);
Signal SumNode_Float232Output_1050: float (5 downto -14);
Signal ProductNode_Float818Output_1051: float (5 downto -14);
Signal ProductNode_Float819weight : float ( 5 downto -14 ) := to_float (0.919660,5,14);

Signal ProductNode_Float819Output_1052: float (5 downto -14);
Signal ProductNode_Float820weight : float ( 5 downto -14 ) := to_float (0.806938,5,14);

Signal ProductNode_Float820Output_1053: float (5 downto -14);
Signal SumNode_Float233Output_1054: float (5 downto -14);
Signal ProductNode_Float821Output_1055: float (5 downto -14);
Signal ProductNode_Float822weight : float ( 5 downto -14 ) := to_float (0.860235,5,14);

Signal ProductNode_Float822Output_1056: float (5 downto -14);
Signal ProductNode_Float823weight : float ( 5 downto -14 ) := to_float (0.941870,5,14);

Signal ProductNode_Float823Output_1057: float (5 downto -14);
Signal ProductNode_Float824weight : float ( 5 downto -14 ) := to_float (0.763101,5,14);

Signal ProductNode_Float824Output_1058: float (5 downto -14);
Signal SumNode_Float234Output_1059: float (5 downto -14);
Signal ProductNode_Float825Output_1060: float (5 downto -14);
Signal SumNode_Float235Output_1061: float (5 downto -14);
Signal ProductNode_Float826Output_1062: float (5 downto -14);
Signal ProductNode_Float827weight : float ( 5 downto -14 ) := to_float (0.693688,5,14);

Signal ProductNode_Float827Output_1063: float (5 downto -14);
Signal ProductNode_Float828weight : float ( 5 downto -14 ) := to_float (0.793165,5,14);

Signal ProductNode_Float828Output_1064: float (5 downto -14);
Signal ProductNode_Float829weight : float ( 5 downto -14 ) := to_float (0.927417,5,14);

Signal ProductNode_Float829Output_1065: float (5 downto -14);
Signal SumNode_Float236Output_1066: float (5 downto -14);
Signal ProductNode_Float830Output_1067: float (5 downto -14);
Signal ProductNode_Float831weight : float ( 5 downto -14 ) := to_float (0.726095,5,14);

Signal ProductNode_Float831Output_1068: float (5 downto -14);
Signal ProductNode_Float832weight : float ( 5 downto -14 ) := to_float (0.909585,5,14);

Signal ProductNode_Float832Output_1069: float (5 downto -14);
Signal ProductNode_Float833weight : float ( 5 downto -14 ) := to_float (0.822920,5,14);

Signal ProductNode_Float833Output_1070: float (5 downto -14);
Signal SumNode_Float237Output_1071: float (5 downto -14);
Signal ProductNode_Float834Output_1072: float (5 downto -14);
Signal ProductNode_Float835weight : float ( 5 downto -14 ) := to_float (0.649155,5,14);

Signal ProductNode_Float835Output_1073: float (5 downto -14);
Signal ProductNode_Float836weight : float ( 5 downto -14 ) := to_float (0.975801,5,14);

Signal ProductNode_Float836Output_1074: float (5 downto -14);
Signal SumNode_Float238Output_1075: float (5 downto -14);
Signal ProductNode_Float837Output_1076: float (5 downto -14);
Signal ProductNode_Float838weight : float ( 5 downto -14 ) := to_float (0.955917,5,14);

Signal ProductNode_Float838Output_1077: float (5 downto -14);
Signal ProductNode_Float839weight : float ( 5 downto -14 ) := to_float (0.790147,5,14);

Signal ProductNode_Float839Output_1078: float (5 downto -14);
Signal ProductNode_Float840weight : float ( 5 downto -14 ) := to_float (0.929014,5,14);

Signal ProductNode_Float840Output_1079: float (5 downto -14);
Signal SumNode_Float239Output_1080: float (5 downto -14);
Signal ProductNode_Float841Output_1081: float (5 downto -14);
Signal SumNode_Float240Output_1082: float (5 downto -14);
Signal ProductNode_Float842Output_1083: float (5 downto -14);
Signal ProductNode_Float843weight : float ( 5 downto -14 ) := to_float (0.965586,5,14);

Signal ProductNode_Float843Output_1084: float (5 downto -14);
Signal SumNode_Float241Output_1085: float (5 downto -14);
Signal ProductNode_Float844Output_1086: float (5 downto -14);
Signal ProductNode_Float845weight : float ( 5 downto -14 ) := to_float (0.750079,5,14);

Signal ProductNode_Float845Output_1087: float (5 downto -14);
Signal ProductNode_Float846weight : float ( 5 downto -14 ) := to_float (0.947231,5,14);

Signal ProductNode_Float846Output_1088: float (5 downto -14);
Signal SumNode_Float242Output_1089: float (5 downto -14);
Signal ProductNode_Float847Output_1090: float (5 downto -14);
Signal ProductNode_Float848weight : float ( 5 downto -14 ) := to_float (0.807766,5,14);

Signal ProductNode_Float848Output_1091: float (5 downto -14);
Signal ProductNode_Float849weight : float ( 5 downto -14 ) := to_float (0.825885,5,14);

Signal ProductNode_Float849Output_1092: float (5 downto -14);
Signal ProductNode_Float850weight : float ( 5 downto -14 ) := to_float (0.617466,5,14);

Signal ProductNode_Float850Output_1093: float (5 downto -14);
Signal ProductNode_Float851weight : float ( 5 downto -14 ) := to_float (0.981367,5,14);

Signal ProductNode_Float851Output_1094: float (5 downto -14);
Signal SumNode_Float243Output_1095: float (5 downto -14);
Signal ProductNode_Float852Output_1096: float (5 downto -14);
Signal ProductNode_Float853weight : float ( 5 downto -14 ) := to_float (0.919167,5,14);

Signal ProductNode_Float853Output_1097: float (5 downto -14);
Signal ProductNode_Float854weight : float ( 5 downto -14 ) := to_float (0.933580,5,14);

Signal ProductNode_Float854Output_1098: float (5 downto -14);
Signal SumNode_Float244Output_1099: float (5 downto -14);
Signal ProductNode_Float855Output_1100: float (5 downto -14);
Signal SumNode_Float245Output_1101: float (5 downto -14);
Signal ProductNode_Float856Output_1102: float (5 downto -14);
Signal ProductNode_Float857weight : float ( 5 downto -14 ) := to_float (0.568305,5,14);

Signal ProductNode_Float857Output_1103: float (5 downto -14);
Signal SumNode_Float246Output_1104: float (5 downto -14);
Signal ProductNode_Float858Output_1105: float (5 downto -14);
Signal ProductNode_Float859weight : float ( 5 downto -14 ) := to_float (0.848299,5,14);

Signal ProductNode_Float859Output_1106: float (5 downto -14);
Signal ProductNode_Float860weight : float ( 5 downto -14 ) := to_float (0.895308,5,14);

Signal ProductNode_Float860Output_1107: float (5 downto -14);
Signal ProductNode_Float861weight : float ( 5 downto -14 ) := to_float (0.842608,5,14);

Signal ProductNode_Float861Output_1108: float (5 downto -14);
Signal SumNode_Float247Output_1109: float (5 downto -14);
Signal ProductNode_Float862Output_1110: float (5 downto -14);
Signal ProductNode_Float863weight : float ( 5 downto -14 ) := to_float (0.870697,5,14);

Signal ProductNode_Float863Output_1111: float (5 downto -14);
Signal ProductNode_Float864weight : float ( 5 downto -14 ) := to_float (0.945793,5,14);

Signal ProductNode_Float864Output_1112: float (5 downto -14);
Signal ProductNode_Float865weight : float ( 5 downto -14 ) := to_float (0.954870,5,14);

Signal ProductNode_Float865Output_1113: float (5 downto -14);
Signal ProductNode_Float866weight : float ( 5 downto -14 ) := to_float (0.870404,5,14);

Signal ProductNode_Float866Output_1114: float (5 downto -14);
Signal ProductNode_Float867weight : float ( 5 downto -14 ) := to_float (0.780732,5,14);

Signal ProductNode_Float867Output_1115: float (5 downto -14);
Signal ProductNode_Float868weight : float ( 5 downto -14 ) := to_float (0.810846,5,14);

Signal ProductNode_Float868Output_1116: float (5 downto -14);
Signal SumNode_Float248Output_1117: float (5 downto -14);
Signal ProductNode_Float869Output_1118: float (5 downto -14);
Signal ProductNode_Float870weight : float ( 5 downto -14 ) := to_float (0.531606,5,14);

Signal ProductNode_Float870Output_1119: float (5 downto -14);
Signal ProductNode_Float871weight : float ( 5 downto -14 ) := to_float (0.669241,5,14);

Signal ProductNode_Float871Output_1120: float (5 downto -14);
Signal ProductNode_Float872weight : float ( 5 downto -14 ) := to_float (0.971580,5,14);

Signal ProductNode_Float872Output_1121: float (5 downto -14);
Signal SumNode_Float249Output_1122: float (5 downto -14);
Signal ProductNode_Float873Output_1123: float (5 downto -14);
Signal ProductNode_Float874weight : float ( 5 downto -14 ) := to_float (0.870697,5,14);

Signal ProductNode_Float874Output_1124: float (5 downto -14);
Signal ProductNode_Float875weight : float ( 5 downto -14 ) := to_float (0.753690,5,14);

Signal ProductNode_Float875Output_1125: float (5 downto -14);
Signal ProductNode_Float876weight : float ( 5 downto -14 ) := to_float (0.774480,5,14);

Signal ProductNode_Float876Output_1126: float (5 downto -14);
Signal ProductNode_Float877weight : float ( 5 downto -14 ) := to_float (0.870404,5,14);

Signal ProductNode_Float877Output_1127: float (5 downto -14);
Signal ProductNode_Float878weight : float ( 5 downto -14 ) := to_float (0.933776,5,14);

Signal ProductNode_Float878Output_1128: float (5 downto -14);
Signal ProductNode_Float879weight : float ( 5 downto -14 ) := to_float (0.660973,5,14);

Signal ProductNode_Float879Output_1129: float (5 downto -14);
Signal SumNode_Float250Output_1130: float (5 downto -14);
Signal ProductNode_Float880Output_1131: float (5 downto -14);
Signal ProductNode_Float881weight : float ( 5 downto -14 ) := to_float (0.870862,5,14);

Signal ProductNode_Float881Output_1132: float (5 downto -14);
Signal SumNode_Float251Output_1133: float (5 downto -14);
Signal ProductNode_Float882Output_1134: float (5 downto -14);
Signal ProductNode_Float883weight : float ( 5 downto -14 ) := to_float (0.888715,5,14);

Signal ProductNode_Float883Output_1135: float (5 downto -14);
Signal ProductNode_Float884weight : float ( 5 downto -14 ) := to_float (0.890735,5,14);

Signal ProductNode_Float884Output_1136: float (5 downto -14);
Signal ProductNode_Float885weight : float ( 5 downto -14 ) := to_float (0.689002,5,14);

Signal ProductNode_Float885Output_1137: float (5 downto -14);
Signal ProductNode_Float886weight : float ( 5 downto -14 ) := to_float (0.966814,5,14);

Signal ProductNode_Float886Output_1138: float (5 downto -14);
Signal SumNode_Float252Output_1139: float (5 downto -14);
Signal ProductNode_Float887Output_1140: float (5 downto -14);
Signal ProductNode_Float888weight : float ( 5 downto -14 ) := to_float (0.551341,5,14);

Signal ProductNode_Float888Output_1141: float (5 downto -14);
Signal ProductNode_Float889weight : float ( 5 downto -14 ) := to_float (0.795357,5,14);

Signal ProductNode_Float889Output_1142: float (5 downto -14);
Signal ProductNode_Float890weight : float ( 5 downto -14 ) := to_float (0.746308,5,14);

Signal ProductNode_Float890Output_1143: float (5 downto -14);
Signal ProductNode_Float891weight : float ( 5 downto -14 ) := to_float (0.989597,5,14);

Signal ProductNode_Float891Output_1144: float (5 downto -14);
Signal ProductNode_Float892weight : float ( 5 downto -14 ) := to_float (0.577708,5,14);

Signal ProductNode_Float892Output_1145: float (5 downto -14);
Signal ProductNode_Float893weight : float ( 5 downto -14 ) := to_float (0.618274,5,14);

Signal ProductNode_Float893Output_1146: float (5 downto -14);
Signal SumNode_Float253Output_1147: float (5 downto -14);
Signal ProductNode_Float894Output_1148: float (5 downto -14);
Signal ProductNode_Float895weight : float ( 5 downto -14 ) := to_float (0.735141,5,14);

Signal ProductNode_Float895Output_1149: float (5 downto -14);
Signal ProductNode_Float896weight : float ( 5 downto -14 ) := to_float (0.495915,5,14);

Signal ProductNode_Float896Output_1150: float (5 downto -14);
Signal ProductNode_Float897weight : float ( 5 downto -14 ) := to_float (0.993928,5,14);

Signal ProductNode_Float897Output_1151: float (5 downto -14);
Signal SumNode_Float254Output_1152: float (5 downto -14);
Signal ProductNode_Float898Output_1153: float (5 downto -14);
Signal ProductNode_Float899weight : float ( 5 downto -14 ) := to_float (0.551341,5,14);

Signal ProductNode_Float899Output_1154: float (5 downto -14);
Signal ProductNode_Float900weight : float ( 5 downto -14 ) := to_float (0.926235,5,14);

Signal ProductNode_Float900Output_1155: float (5 downto -14);
Signal ProductNode_Float901weight : float ( 5 downto -14 ) := to_float (0.616494,5,14);

Signal ProductNode_Float901Output_1156: float (5 downto -14);
Signal ProductNode_Float902weight : float ( 5 downto -14 ) := to_float (0.989597,5,14);

Signal ProductNode_Float902Output_1157: float (5 downto -14);
Signal ProductNode_Float903weight : float ( 5 downto -14 ) := to_float (0.986786,5,14);

Signal ProductNode_Float903Output_1158: float (5 downto -14);
Signal ProductNode_Float904weight : float ( 5 downto -14 ) := to_float (0.464416,5,14);

Signal ProductNode_Float904Output_1159: float (5 downto -14);
Signal SumNode_Float255Output_1160: float (5 downto -14);
Signal ProductNode_Float905Output_1161: float (5 downto -14);
Signal ProductNode_Float906weight : float ( 5 downto -14 ) := to_float (0.938375,5,14);

Signal ProductNode_Float906Output_1162: float (5 downto -14);
Signal SumNode_Float256Output_1163: float (5 downto -14);
Signal ProductNode_Float907Output_1164: float (5 downto -14);
Signal ProductNode_Float908weight : float ( 5 downto -14 ) := to_float (0.978422,5,14);

Signal ProductNode_Float908Output_1165: float (5 downto -14);
Signal SumNode_Float257Output_1166: float (5 downto -14);
Signal ProductNode_Float909Output_1167: float (5 downto -14);
Signal ProductNode_Float910weight : float ( 5 downto -14 ) := to_float (0.773183,5,14);

Signal ProductNode_Float910Output_1168: float (5 downto -14);
Signal ProductNode_Float911weight : float ( 5 downto -14 ) := to_float (0.848299,5,14);

Signal ProductNode_Float911Output_1169: float (5 downto -14);
Signal ProductNode_Float912weight : float ( 5 downto -14 ) := to_float (0.562709,5,14);

Signal ProductNode_Float912Output_1170: float (5 downto -14);
Signal ProductNode_Float913weight : float ( 5 downto -14 ) := to_float (0.988453,5,14);

Signal ProductNode_Float913Output_1171: float (5 downto -14);
Signal SumNode_Float258Output_1172: float (5 downto -14);
Signal ProductNode_Float914Output_1173: float (5 downto -14);
Signal ProductNode_Float915weight : float ( 5 downto -14 ) := to_float (0.870697,5,14);

Signal ProductNode_Float915Output_1174: float (5 downto -14);
Signal ProductNode_Float916weight : float ( 5 downto -14 ) := to_float (0.945793,5,14);

Signal ProductNode_Float916Output_1175: float (5 downto -14);
Signal ProductNode_Float917weight : float ( 5 downto -14 ) := to_float (0.729204,5,14);

Signal ProductNode_Float917Output_1176: float (5 downto -14);
Signal ProductNode_Float918weight : float ( 5 downto -14 ) := to_float (0.870404,5,14);

Signal ProductNode_Float918Output_1177: float (5 downto -14);
Signal ProductNode_Float919weight : float ( 5 downto -14 ) := to_float (0.780732,5,14);

Signal ProductNode_Float919Output_1178: float (5 downto -14);
Signal ProductNode_Float920weight : float ( 5 downto -14 ) := to_float (0.917308,5,14);

Signal ProductNode_Float920Output_1179: float (5 downto -14);
Signal SumNode_Float259Output_1180: float (5 downto -14);
Signal ProductNode_Float921Output_1181: float (5 downto -14);
Signal ProductNode_Float922weight : float ( 5 downto -14 ) := to_float (0.631626,5,14);

Signal ProductNode_Float922Output_1182: float (5 downto -14);
Signal ProductNode_Float923weight : float ( 5 downto -14 ) := to_float (0.453222,5,14);

Signal ProductNode_Float923Output_1183: float (5 downto -14);
Signal ProductNode_Float924weight : float ( 5 downto -14 ) := to_float (0.996146,5,14);

Signal ProductNode_Float924Output_1184: float (5 downto -14);
Signal SumNode_Float260Output_1185: float (5 downto -14);
Signal ProductNode_Float925Output_1186: float (5 downto -14);
Signal ProductNode_Float926weight : float ( 5 downto -14 ) := to_float (0.870697,5,14);

Signal ProductNode_Float926Output_1187: float (5 downto -14);
Signal ProductNode_Float927weight : float ( 5 downto -14 ) := to_float (0.753690,5,14);

Signal ProductNode_Float927Output_1188: float (5 downto -14);
Signal ProductNode_Float928weight : float ( 5 downto -14 ) := to_float (0.936763,5,14);

Signal ProductNode_Float928Output_1189: float (5 downto -14);
Signal ProductNode_Float929weight : float ( 5 downto -14 ) := to_float (0.870404,5,14);

Signal ProductNode_Float929Output_1190: float (5 downto -14);
Signal ProductNode_Float930weight : float ( 5 downto -14 ) := to_float (0.933776,5,14);

Signal ProductNode_Float930Output_1191: float (5 downto -14);
Signal ProductNode_Float931weight : float ( 5 downto -14 ) := to_float (0.973389,5,14);

Signal ProductNode_Float931Output_1192: float (5 downto -14);
Signal SumNode_Float261Output_1193: float (5 downto -14);
Signal ProductNode_Float932Output_1194: float (5 downto -14);
Signal ProductNode_Float933weight : float ( 5 downto -14 ) := to_float (0.912549,5,14);

Signal ProductNode_Float933Output_1195: float (5 downto -14);
Signal SumNode_Float262Output_1196: float (5 downto -14);
Signal ProductNode_Float934Output_1197: float (5 downto -14);
Signal ProductNode_Float935weight : float ( 5 downto -14 ) := to_float (0.973991,5,14);

Signal ProductNode_Float935Output_1198: float (5 downto -14);
Signal ProductNode_Float936weight : float ( 5 downto -14 ) := to_float (0.890735,5,14);

Signal ProductNode_Float936Output_1199: float (5 downto -14);
Signal ProductNode_Float937weight : float ( 5 downto -14 ) := to_float (0.382644,5,14);

Signal ProductNode_Float937Output_1200: float (5 downto -14);
Signal ProductNode_Float938weight : float ( 5 downto -14 ) := to_float (0.998354,5,14);

Signal ProductNode_Float938Output_1201: float (5 downto -14);
Signal SumNode_Float263Output_1202: float (5 downto -14);
Signal ProductNode_Float939Output_1203: float (5 downto -14);
Signal ProductNode_Float940weight : float ( 5 downto -14 ) := to_float (0.551341,5,14);

Signal ProductNode_Float940Output_1204: float (5 downto -14);
Signal ProductNode_Float941weight : float ( 5 downto -14 ) := to_float (0.795357,5,14);

Signal ProductNode_Float941Output_1205: float (5 downto -14);
Signal ProductNode_Float942weight : float ( 5 downto -14 ) := to_float (0.948695,5,14);

Signal ProductNode_Float942Output_1206: float (5 downto -14);
Signal ProductNode_Float943weight : float ( 5 downto -14 ) := to_float (0.989597,5,14);

Signal ProductNode_Float943Output_1207: float (5 downto -14);
Signal ProductNode_Float944weight : float ( 5 downto -14 ) := to_float (0.577708,5,14);

Signal ProductNode_Float944Output_1208: float (5 downto -14);
Signal ProductNode_Float945weight : float ( 5 downto -14 ) := to_float (0.981240,5,14);

Signal ProductNode_Float945Output_1209: float (5 downto -14);
Signal SumNode_Float264Output_1210: float (5 downto -14);
Signal ProductNode_Float946Output_1211: float (5 downto -14);
Signal ProductNode_Float947weight : float ( 5 downto -14 ) := to_float (0.712179,5,14);

Signal ProductNode_Float947Output_1212: float (5 downto -14);
Signal ProductNode_Float948weight : float ( 5 downto -14 ) := to_float (0.336149,5,14);

Signal ProductNode_Float948Output_1213: float (5 downto -14);
Signal ProductNode_Float949weight : float ( 5 downto -14 ) := to_float (0.999140,5,14);

Signal ProductNode_Float949Output_1214: float (5 downto -14);
Signal SumNode_Float265Output_1215: float (5 downto -14);
Signal ProductNode_Float950Output_1216: float (5 downto -14);
Signal ProductNode_Float951weight : float ( 5 downto -14 ) := to_float (0.551341,5,14);

Signal ProductNode_Float951Output_1217: float (5 downto -14);
Signal ProductNode_Float952weight : float ( 5 downto -14 ) := to_float (0.926235,5,14);

Signal ProductNode_Float952Output_1218: float (5 downto -14);
Signal ProductNode_Float953weight : float ( 5 downto -14 ) := to_float (0.981519,5,14);

Signal ProductNode_Float953Output_1219: float (5 downto -14);
Signal ProductNode_Float954weight : float ( 5 downto -14 ) := to_float (0.989597,5,14);

Signal ProductNode_Float954Output_1220: float (5 downto -14);
Signal ProductNode_Float955weight : float ( 5 downto -14 ) := to_float (0.986786,5,14);

Signal ProductNode_Float955Output_1221: float (5 downto -14);
Signal ProductNode_Float956weight : float ( 5 downto -14 ) := to_float (0.995641,5,14);

Signal ProductNode_Float956Output_1222: float (5 downto -14);
Signal SumNode_Float266Output_1223: float (5 downto -14);
Signal ProductNode_Float957Output_1224: float (5 downto -14);
Signal ProductNode_Float958weight : float ( 5 downto -14 ) := to_float (0.972670,5,14);

Signal ProductNode_Float958Output_1225: float (5 downto -14);
Signal SumNode_Float267Output_1226: float (5 downto -14);
Signal ProductNode_Float959Output_1227: float (5 downto -14);
Signal ProductNode_Float960weight : float ( 5 downto -14 ) := to_float (0.991382,5,14);

Signal ProductNode_Float960Output_1228: float (5 downto -14);
Signal SumNode_Float268Output_1229: float (5 downto -14);
Signal ProductNode_Float961Output_1230: float (5 downto -14);
Signal ProductNode_Float962weight : float ( 5 downto -14 ) := to_float (0.569080,5,14);

Signal ProductNode_Float962Output_1231: float (5 downto -14);
Signal SumNode_Float269Output_1232: float (5 downto -14);
Signal ProductNode_Float963Output_1233: float (5 downto -14);
Signal ProductNode_Float964weight : float ( 5 downto -14 ) := to_float (0.965849,5,14);

Signal ProductNode_Float964Output_1234: float (5 downto -14);
Signal ProductNode_Float965weight : float ( 5 downto -14 ) := to_float (0.692695,5,14);

Signal ProductNode_Float965Output_1235: float (5 downto -14);
Signal SumNode_Float270Output_1236: float (5 downto -14);
Signal ProductNode_Float966Output_1237: float (5 downto -14);
Signal ProductNode_Float967weight : float ( 5 downto -14 ) := to_float (0.880399,5,14);

Signal ProductNode_Float967Output_1238: float (5 downto -14);
Signal ProductNode_Float968weight : float ( 5 downto -14 ) := to_float (0.997554,5,14);

Signal ProductNode_Float968Output_1239: float (5 downto -14);
Signal ProductNode_Float969weight : float ( 5 downto -14 ) := to_float (0.414069,5,14);

Signal ProductNode_Float969Output_1240: float (5 downto -14);
Signal SumNode_Float271Output_1241: float (5 downto -14);
Signal ProductNode_Float970Output_1242: float (5 downto -14);
Signal ProductNode_Float971weight : float ( 5 downto -14 ) := to_float (0.919660,5,14);

Signal ProductNode_Float971Output_1243: float (5 downto -14);
Signal ProductNode_Float972weight : float ( 5 downto -14 ) := to_float (0.806938,5,14);

Signal ProductNode_Float972Output_1244: float (5 downto -14);
Signal SumNode_Float272Output_1245: float (5 downto -14);
Signal ProductNode_Float973Output_1246: float (5 downto -14);
Signal ProductNode_Float974weight : float ( 5 downto -14 ) := to_float (0.860235,5,14);

Signal ProductNode_Float974Output_1247: float (5 downto -14);
Signal ProductNode_Float975weight : float ( 5 downto -14 ) := to_float (0.989739,5,14);

Signal ProductNode_Float975Output_1248: float (5 downto -14);
Signal ProductNode_Float976weight : float ( 5 downto -14 ) := to_float (0.549861,5,14);

Signal ProductNode_Float976Output_1249: float (5 downto -14);
Signal SumNode_Float273Output_1250: float (5 downto -14);
Signal ProductNode_Float977Output_1251: float (5 downto -14);
Signal SumNode_Float274Output_1252: float (5 downto -14);
Signal ProductNode_Float978Output_1253: float (5 downto -14);
Signal ProductNode_Float979weight : float ( 5 downto -14 ) := to_float (0.984104,5,14);

Signal ProductNode_Float979Output_1254: float (5 downto -14);
Signal ProductNode_Float980weight : float ( 5 downto -14 ) := to_float (0.793165,5,14);

Signal ProductNode_Float980Output_1255: float (5 downto -14);
Signal ProductNode_Float981weight : float ( 5 downto -14 ) := to_float (0.927417,5,14);

Signal ProductNode_Float981Output_1256: float (5 downto -14);
Signal SumNode_Float275Output_1257: float (5 downto -14);
Signal ProductNode_Float982Output_1258: float (5 downto -14);
Signal ProductNode_Float983weight : float ( 5 downto -14 ) := to_float (0.726095,5,14);

Signal ProductNode_Float983Output_1259: float (5 downto -14);
Signal ProductNode_Float984weight : float ( 5 downto -14 ) := to_float (0.988880,5,14);

Signal ProductNode_Float984Output_1260: float (5 downto -14);
Signal ProductNode_Float985weight : float ( 5 downto -14 ) := to_float (0.558577,5,14);

Signal ProductNode_Float985Output_1261: float (5 downto -14);
Signal SumNode_Float276Output_1262: float (5 downto -14);
Signal ProductNode_Float986Output_1263: float (5 downto -14);
Signal ProductNode_Float987weight : float ( 5 downto -14 ) := to_float (0.649155,5,14);

Signal ProductNode_Float987Output_1264: float (5 downto -14);
Signal ProductNode_Float988weight : float ( 5 downto -14 ) := to_float (0.975801,5,14);

Signal ProductNode_Float988Output_1265: float (5 downto -14);
Signal SumNode_Float277Output_1266: float (5 downto -14);
Signal ProductNode_Float989Output_1267: float (5 downto -14);
Signal ProductNode_Float990weight : float ( 5 downto -14 ) := to_float (0.955917,5,14);

Signal ProductNode_Float990Output_1268: float (5 downto -14);
Signal ProductNode_Float991weight : float ( 5 downto -14 ) := to_float (0.985013,5,14);

Signal ProductNode_Float991Output_1269: float (5 downto -14);
Signal ProductNode_Float992weight : float ( 5 downto -14 ) := to_float (0.592017,5,14);

Signal ProductNode_Float992Output_1270: float (5 downto -14);
Signal SumNode_Float278Output_1271: float (5 downto -14);
Signal ProductNode_Float993Output_1272: float (5 downto -14);
Signal SumNode_Float279Output_1273: float (5 downto -14);
Signal ProductNode_Float994Output_1274: float (5 downto -14);
Signal ProductNode_Float995weight : float ( 5 downto -14 ) := to_float (0.598812,5,14);

Signal ProductNode_Float995Output_1275: float (5 downto -14);
Signal SumNode_Float280Output_1276: float (5 downto -14);
Signal ProductNode_Float996Output_1277: float (5 downto -14);
Signal ProductNode_Float997weight : float ( 5 downto -14 ) := to_float (0.927615,5,14);

Signal ProductNode_Float997Output_1278: float (5 downto -14);
Signal ProductNode_Float998weight : float ( 5 downto -14 ) := to_float (0.792795,5,14);

Signal ProductNode_Float998Output_1279: float (5 downto -14);
Signal SumNode_Float281Output_1280: float (5 downto -14);
Signal ProductNode_Float999Output_1281: float (5 downto -14);
Signal ProductNode_Float1000weight : float ( 5 downto -14 ) := to_float (0.907425,5,14);

Signal ProductNode_Float1000Output_1282: float (5 downto -14);
Signal ProductNode_Float1001weight : float ( 5 downto -14 ) := to_float (0.948402,5,14);

Signal ProductNode_Float1001Output_1283: float (5 downto -14);
Signal ProductNode_Float1002weight : float ( 5 downto -14 ) := to_float (0.838940,5,14);

Signal ProductNode_Float1002Output_1284: float (5 downto -14);
Signal ProductNode_Float1003weight : float ( 5 downto -14 ) := to_float (0.898142,5,14);

Signal ProductNode_Float1003Output_1285: float (5 downto -14);
Signal SumNode_Float282Output_1286: float (5 downto -14);
Signal ProductNode_Float1004Output_1287: float (5 downto -14);
Signal ProductNode_Float1005weight : float ( 5 downto -14 ) := to_float (0.826105,5,14);

Signal ProductNode_Float1005Output_1288: float (5 downto -14);
Signal ProductNode_Float1006weight : float ( 5 downto -14 ) := to_float (0.838083,5,14);

Signal ProductNode_Float1006Output_1289: float (5 downto -14);
Signal SumNode_Float283Output_1290: float (5 downto -14);
Signal ProductNode_Float1007Output_1291: float (5 downto -14);
Signal ProductNode_Float1008weight : float ( 5 downto -14 ) := to_float (0.965849,5,14);

Signal ProductNode_Float1008Output_1292: float (5 downto -14);
Signal ProductNode_Float1009weight : float ( 5 downto -14 ) := to_float (0.692695,5,14);

Signal ProductNode_Float1009Output_1293: float (5 downto -14);
Signal SumNode_Float284Output_1294: float (5 downto -14);
Signal ProductNode_Float1010Output_1295: float (5 downto -14);
Signal ProductNode_Float1011weight : float ( 5 downto -14 ) := to_float (0.880399,5,14);

Signal ProductNode_Float1011Output_1296: float (5 downto -14);
Signal ProductNode_Float1012weight : float ( 5 downto -14 ) := to_float (0.997554,5,14);

Signal ProductNode_Float1012Output_1297: float (5 downto -14);
Signal ProductNode_Float1013weight : float ( 5 downto -14 ) := to_float (0.414069,5,14);

Signal ProductNode_Float1013Output_1298: float (5 downto -14);
Signal SumNode_Float285Output_1299: float (5 downto -14);
Signal ProductNode_Float1014Output_1300: float (5 downto -14);
Signal ProductNode_Float1015weight : float ( 5 downto -14 ) := to_float (0.919660,5,14);

Signal ProductNode_Float1015Output_1301: float (5 downto -14);
Signal ProductNode_Float1016weight : float ( 5 downto -14 ) := to_float (0.806938,5,14);

Signal ProductNode_Float1016Output_1302: float (5 downto -14);
Signal SumNode_Float286Output_1303: float (5 downto -14);
Signal ProductNode_Float1017Output_1304: float (5 downto -14);
Signal ProductNode_Float1018weight : float ( 5 downto -14 ) := to_float (0.860235,5,14);

Signal ProductNode_Float1018Output_1305: float (5 downto -14);
Signal ProductNode_Float1019weight : float ( 5 downto -14 ) := to_float (0.989739,5,14);

Signal ProductNode_Float1019Output_1306: float (5 downto -14);
Signal ProductNode_Float1020weight : float ( 5 downto -14 ) := to_float (0.549861,5,14);

Signal ProductNode_Float1020Output_1307: float (5 downto -14);
Signal SumNode_Float287Output_1308: float (5 downto -14);
Signal ProductNode_Float1021Output_1309: float (5 downto -14);
Signal SumNode_Float288Output_1310: float (5 downto -14);
Signal ProductNode_Float1022Output_1311: float (5 downto -14);
Signal ProductNode_Float1023weight : float ( 5 downto -14 ) := to_float (0.932937,5,14);

Signal ProductNode_Float1023Output_1312: float (5 downto -14);
Signal ProductNode_Float1024weight : float ( 5 downto -14 ) := to_float (0.793165,5,14);

Signal ProductNode_Float1024Output_1313: float (5 downto -14);
Signal ProductNode_Float1025weight : float ( 5 downto -14 ) := to_float (0.927417,5,14);

Signal ProductNode_Float1025Output_1314: float (5 downto -14);
Signal SumNode_Float289Output_1315: float (5 downto -14);
Signal ProductNode_Float1026Output_1316: float (5 downto -14);
Signal ProductNode_Float1027weight : float ( 5 downto -14 ) := to_float (0.726095,5,14);

Signal ProductNode_Float1027Output_1317: float (5 downto -14);
Signal ProductNode_Float1028weight : float ( 5 downto -14 ) := to_float (0.988880,5,14);

Signal ProductNode_Float1028Output_1318: float (5 downto -14);
Signal ProductNode_Float1029weight : float ( 5 downto -14 ) := to_float (0.558577,5,14);

Signal ProductNode_Float1029Output_1319: float (5 downto -14);
Signal SumNode_Float290Output_1320: float (5 downto -14);
Signal ProductNode_Float1030Output_1321: float (5 downto -14);
Signal ProductNode_Float1031weight : float ( 5 downto -14 ) := to_float (0.649155,5,14);

Signal ProductNode_Float1031Output_1322: float (5 downto -14);
Signal ProductNode_Float1032weight : float ( 5 downto -14 ) := to_float (0.975801,5,14);

Signal ProductNode_Float1032Output_1323: float (5 downto -14);
Signal SumNode_Float291Output_1324: float (5 downto -14);
Signal ProductNode_Float1033Output_1325: float (5 downto -14);
Signal ProductNode_Float1034weight : float ( 5 downto -14 ) := to_float (0.955917,5,14);

Signal ProductNode_Float1034Output_1326: float (5 downto -14);
Signal ProductNode_Float1035weight : float ( 5 downto -14 ) := to_float (0.985013,5,14);

Signal ProductNode_Float1035Output_1327: float (5 downto -14);
Signal ProductNode_Float1036weight : float ( 5 downto -14 ) := to_float (0.592017,5,14);

Signal ProductNode_Float1036Output_1328: float (5 downto -14);
Signal SumNode_Float292Output_1329: float (5 downto -14);
Signal ProductNode_Float1037Output_1330: float (5 downto -14);
Signal SumNode_Float293Output_1331: float (5 downto -14);
Signal ProductNode_Float1038Output_1332: float (5 downto -14);
Signal ProductNode_Float1039weight : float ( 5 downto -14 ) := to_float (0.782438,5,14);

Signal ProductNode_Float1039Output_1333: float (5 downto -14);
Signal SumNode_Float294Output_1334: float (5 downto -14);
Signal ProductNode_Float1040Output_1335: float (5 downto -14);
Signal ProductNode_Float1041weight : float ( 5 downto -14 ) := to_float (0.750079,5,14);

Signal ProductNode_Float1041Output_1336: float (5 downto -14);
Signal ProductNode_Float1042weight : float ( 5 downto -14 ) := to_float (0.947231,5,14);

Signal ProductNode_Float1042Output_1337: float (5 downto -14);
Signal SumNode_Float295Output_1338: float (5 downto -14);
Signal ProductNode_Float1043Output_1339: float (5 downto -14);
Signal ProductNode_Float1044weight : float ( 5 downto -14 ) := to_float (0.907425,5,14);

Signal ProductNode_Float1044Output_1340: float (5 downto -14);
Signal ProductNode_Float1045weight : float ( 5 downto -14 ) := to_float (0.747070,5,14);

Signal ProductNode_Float1045Output_1341: float (5 downto -14);
Signal ProductNode_Float1046weight : float ( 5 downto -14 ) := to_float (0.617466,5,14);

Signal ProductNode_Float1046Output_1342: float (5 downto -14);
Signal ProductNode_Float1047weight : float ( 5 downto -14 ) := to_float (0.981367,5,14);

Signal ProductNode_Float1047Output_1343: float (5 downto -14);
Signal SumNode_Float296Output_1344: float (5 downto -14);
Signal ProductNode_Float1048Output_1345: float (5 downto -14);
Signal ProductNode_Float1049weight : float ( 5 downto -14 ) := to_float (0.826105,5,14);

Signal ProductNode_Float1049Output_1346: float (5 downto -14);
Signal ProductNode_Float1050weight : float ( 5 downto -14 ) := to_float (0.898792,5,14);

Signal ProductNode_Float1050Output_1347: float (5 downto -14);
Signal SumNode_Float297Output_1348: float (5 downto -14);
Signal ProductNode_Float1051Output_1349: float (5 downto -14);
Signal SumNode_Float298Output_1350: float (5 downto -14);
Signal ProductNode_Float1052Output_1351: float (5 downto -14);
Signal ProductNode_Float1053weight : float ( 5 downto -14 ) := to_float (0.914453,5,14);

Signal ProductNode_Float1053Output_1352: float (5 downto -14);
Signal ProductNode_Float1054weight : float ( 5 downto -14 ) := to_float (0.965849,5,14);

Signal ProductNode_Float1054Output_1353: float (5 downto -14);
Signal ProductNode_Float1055weight : float ( 5 downto -14 ) := to_float (0.692695,5,14);

Signal ProductNode_Float1055Output_1354: float (5 downto -14);
Signal SumNode_Float299Output_1355: float (5 downto -14);
Signal ProductNode_Float1056Output_1356: float (5 downto -14);
Signal ProductNode_Float1057weight : float ( 5 downto -14 ) := to_float (0.880399,5,14);

Signal ProductNode_Float1057Output_1357: float (5 downto -14);
Signal ProductNode_Float1058weight : float ( 5 downto -14 ) := to_float (0.966381,5,14);

Signal ProductNode_Float1058Output_1358: float (5 downto -14);
Signal ProductNode_Float1059weight : float ( 5 downto -14 ) := to_float (0.690672,5,14);

Signal ProductNode_Float1059Output_1359: float (5 downto -14);
Signal SumNode_Float300Output_1360: float (5 downto -14);
Signal ProductNode_Float1060Output_1361: float (5 downto -14);
Signal ProductNode_Float1061weight : float ( 5 downto -14 ) := to_float (0.919660,5,14);

Signal ProductNode_Float1061Output_1362: float (5 downto -14);
Signal ProductNode_Float1062weight : float ( 5 downto -14 ) := to_float (0.806938,5,14);

Signal ProductNode_Float1062Output_1363: float (5 downto -14);
Signal SumNode_Float301Output_1364: float (5 downto -14);
Signal ProductNode_Float1063Output_1365: float (5 downto -14);
Signal ProductNode_Float1064weight : float ( 5 downto -14 ) := to_float (0.860235,5,14);

Signal ProductNode_Float1064Output_1366: float (5 downto -14);
Signal ProductNode_Float1065weight : float ( 5 downto -14 ) := to_float (0.941870,5,14);

Signal ProductNode_Float1065Output_1367: float (5 downto -14);
Signal ProductNode_Float1066weight : float ( 5 downto -14 ) := to_float (0.763101,5,14);

Signal ProductNode_Float1066Output_1368: float (5 downto -14);
Signal SumNode_Float302Output_1369: float (5 downto -14);
Signal ProductNode_Float1067Output_1370: float (5 downto -14);
Signal SumNode_Float303Output_1371: float (5 downto -14);
Signal ProductNode_Float1068Output_1372: float (5 downto -14);
Signal ProductNode_Float1069weight : float ( 5 downto -14 ) := to_float (0.924413,5,14);

Signal ProductNode_Float1069Output_1373: float (5 downto -14);
Signal ProductNode_Float1070weight : float ( 5 downto -14 ) := to_float (0.793165,5,14);

Signal ProductNode_Float1070Output_1374: float (5 downto -14);
Signal ProductNode_Float1071weight : float ( 5 downto -14 ) := to_float (0.927417,5,14);

Signal ProductNode_Float1071Output_1375: float (5 downto -14);
Signal SumNode_Float304Output_1376: float (5 downto -14);
Signal ProductNode_Float1072Output_1377: float (5 downto -14);
Signal ProductNode_Float1073weight : float ( 5 downto -14 ) := to_float (0.726095,5,14);

Signal ProductNode_Float1073Output_1378: float (5 downto -14);
Signal ProductNode_Float1074weight : float ( 5 downto -14 ) := to_float (0.909585,5,14);

Signal ProductNode_Float1074Output_1379: float (5 downto -14);
Signal ProductNode_Float1075weight : float ( 5 downto -14 ) := to_float (0.822920,5,14);

Signal ProductNode_Float1075Output_1380: float (5 downto -14);
Signal SumNode_Float305Output_1381: float (5 downto -14);
Signal ProductNode_Float1076Output_1382: float (5 downto -14);
Signal ProductNode_Float1077weight : float ( 5 downto -14 ) := to_float (0.649155,5,14);

Signal ProductNode_Float1077Output_1383: float (5 downto -14);
Signal ProductNode_Float1078weight : float ( 5 downto -14 ) := to_float (0.975801,5,14);

Signal ProductNode_Float1078Output_1384: float (5 downto -14);
Signal SumNode_Float306Output_1385: float (5 downto -14);
Signal ProductNode_Float1079Output_1386: float (5 downto -14);
Signal ProductNode_Float1080weight : float ( 5 downto -14 ) := to_float (0.955917,5,14);

Signal ProductNode_Float1080Output_1387: float (5 downto -14);
Signal ProductNode_Float1081weight : float ( 5 downto -14 ) := to_float (0.790147,5,14);

Signal ProductNode_Float1081Output_1388: float (5 downto -14);
Signal ProductNode_Float1082weight : float ( 5 downto -14 ) := to_float (0.929014,5,14);

Signal ProductNode_Float1082Output_1389: float (5 downto -14);
Signal SumNode_Float307Output_1390: float (5 downto -14);
Signal ProductNode_Float1083Output_1391: float (5 downto -14);
Signal SumNode_Float308Output_1392: float (5 downto -14);
Signal ProductNode_Float1084Output_1393: float (5 downto -14);
Signal ProductNode_Float1085weight : float ( 5 downto -14 ) := to_float (0.798666,5,14);

Signal ProductNode_Float1085Output_1394: float (5 downto -14);
Signal SumNode_Float309Output_1395: float (5 downto -14);
Signal ProductNode_Float1086Output_1396: float (5 downto -14);
Signal ProductNode_Float1087weight : float ( 5 downto -14 ) := to_float (0.927615,5,14);

Signal ProductNode_Float1087Output_1397: float (5 downto -14);
Signal ProductNode_Float1088weight : float ( 5 downto -14 ) := to_float (0.792795,5,14);

Signal ProductNode_Float1088Output_1398: float (5 downto -14);
Signal SumNode_Float310Output_1399: float (5 downto -14);
Signal ProductNode_Float1089Output_1400: float (5 downto -14);
Signal ProductNode_Float1090weight : float ( 5 downto -14 ) := to_float (0.807766,5,14);

Signal ProductNode_Float1090Output_1401: float (5 downto -14);
Signal ProductNode_Float1091weight : float ( 5 downto -14 ) := to_float (0.907576,5,14);

Signal ProductNode_Float1091Output_1402: float (5 downto -14);
Signal ProductNode_Float1092weight : float ( 5 downto -14 ) := to_float (0.838940,5,14);

Signal ProductNode_Float1092Output_1403: float (5 downto -14);
Signal ProductNode_Float1093weight : float ( 5 downto -14 ) := to_float (0.898142,5,14);

Signal ProductNode_Float1093Output_1404: float (5 downto -14);
Signal SumNode_Float311Output_1405: float (5 downto -14);
Signal ProductNode_Float1094Output_1406: float (5 downto -14);
Signal ProductNode_Float1095weight : float ( 5 downto -14 ) := to_float (0.919167,5,14);

Signal ProductNode_Float1095Output_1407: float (5 downto -14);
Signal ProductNode_Float1096weight : float ( 5 downto -14 ) := to_float (0.781132,5,14);

Signal ProductNode_Float1096Output_1408: float (5 downto -14);
Signal SumNode_Float312Output_1409: float (5 downto -14);
Signal ProductNode_Float1097Output_1410: float (5 downto -14);
Signal ProductNode_Float1098weight : float ( 5 downto -14 ) := to_float (0.965849,5,14);

Signal ProductNode_Float1098Output_1411: float (5 downto -14);
Signal ProductNode_Float1099weight : float ( 5 downto -14 ) := to_float (0.692695,5,14);

Signal ProductNode_Float1099Output_1412: float (5 downto -14);
Signal SumNode_Float313Output_1413: float (5 downto -14);
Signal ProductNode_Float1100Output_1414: float (5 downto -14);
Signal ProductNode_Float1101weight : float ( 5 downto -14 ) := to_float (0.880399,5,14);

Signal ProductNode_Float1101Output_1415: float (5 downto -14);
Signal ProductNode_Float1102weight : float ( 5 downto -14 ) := to_float (0.966381,5,14);

Signal ProductNode_Float1102Output_1416: float (5 downto -14);
Signal ProductNode_Float1103weight : float ( 5 downto -14 ) := to_float (0.690672,5,14);

Signal ProductNode_Float1103Output_1417: float (5 downto -14);
Signal SumNode_Float314Output_1418: float (5 downto -14);
Signal ProductNode_Float1104Output_1419: float (5 downto -14);
Signal ProductNode_Float1105weight : float ( 5 downto -14 ) := to_float (0.919660,5,14);

Signal ProductNode_Float1105Output_1420: float (5 downto -14);
Signal ProductNode_Float1106weight : float ( 5 downto -14 ) := to_float (0.806938,5,14);

Signal ProductNode_Float1106Output_1421: float (5 downto -14);
Signal SumNode_Float315Output_1422: float (5 downto -14);
Signal ProductNode_Float1107Output_1423: float (5 downto -14);
Signal ProductNode_Float1108weight : float ( 5 downto -14 ) := to_float (0.860235,5,14);

Signal ProductNode_Float1108Output_1424: float (5 downto -14);
Signal ProductNode_Float1109weight : float ( 5 downto -14 ) := to_float (0.941870,5,14);

Signal ProductNode_Float1109Output_1425: float (5 downto -14);
Signal ProductNode_Float1110weight : float ( 5 downto -14 ) := to_float (0.763101,5,14);

Signal ProductNode_Float1110Output_1426: float (5 downto -14);
Signal SumNode_Float316Output_1427: float (5 downto -14);
Signal ProductNode_Float1111Output_1428: float (5 downto -14);
Signal SumNode_Float317Output_1429: float (5 downto -14);
Signal ProductNode_Float1112Output_1430: float (5 downto -14);
Signal ProductNode_Float1113weight : float ( 5 downto -14 ) := to_float (0.693688,5,14);

Signal ProductNode_Float1113Output_1431: float (5 downto -14);
Signal ProductNode_Float1114weight : float ( 5 downto -14 ) := to_float (0.793165,5,14);

Signal ProductNode_Float1114Output_1432: float (5 downto -14);
Signal ProductNode_Float1115weight : float ( 5 downto -14 ) := to_float (0.927417,5,14);

Signal ProductNode_Float1115Output_1433: float (5 downto -14);
Signal SumNode_Float318Output_1434: float (5 downto -14);
Signal ProductNode_Float1116Output_1435: float (5 downto -14);
Signal ProductNode_Float1117weight : float ( 5 downto -14 ) := to_float (0.726095,5,14);

Signal ProductNode_Float1117Output_1436: float (5 downto -14);
Signal ProductNode_Float1118weight : float ( 5 downto -14 ) := to_float (0.909585,5,14);

Signal ProductNode_Float1118Output_1437: float (5 downto -14);
Signal ProductNode_Float1119weight : float ( 5 downto -14 ) := to_float (0.822920,5,14);

Signal ProductNode_Float1119Output_1438: float (5 downto -14);
Signal SumNode_Float319Output_1439: float (5 downto -14);
Signal ProductNode_Float1120Output_1440: float (5 downto -14);
Signal ProductNode_Float1121weight : float ( 5 downto -14 ) := to_float (0.649155,5,14);

Signal ProductNode_Float1121Output_1441: float (5 downto -14);
Signal ProductNode_Float1122weight : float ( 5 downto -14 ) := to_float (0.975801,5,14);

Signal ProductNode_Float1122Output_1442: float (5 downto -14);
Signal SumNode_Float320Output_1443: float (5 downto -14);
Signal ProductNode_Float1123Output_1444: float (5 downto -14);
Signal ProductNode_Float1124weight : float ( 5 downto -14 ) := to_float (0.955917,5,14);

Signal ProductNode_Float1124Output_1445: float (5 downto -14);
Signal ProductNode_Float1125weight : float ( 5 downto -14 ) := to_float (0.790147,5,14);

Signal ProductNode_Float1125Output_1446: float (5 downto -14);
Signal ProductNode_Float1126weight : float ( 5 downto -14 ) := to_float (0.929014,5,14);

Signal ProductNode_Float1126Output_1447: float (5 downto -14);
Signal SumNode_Float321Output_1448: float (5 downto -14);
Signal ProductNode_Float1127Output_1449: float (5 downto -14);
Signal SumNode_Float322Output_1450: float (5 downto -14);
Signal ProductNode_Float1128Output_1451: float (5 downto -14);
Signal ProductNode_Float1129weight : float ( 5 downto -14 ) := to_float (0.965586,5,14);

Signal ProductNode_Float1129Output_1452: float (5 downto -14);
Signal SumNode_Float323Output_1453: float (5 downto -14);
Signal ProductNode_Float1130Output_1454: float (5 downto -14);
Signal ProductNode_Float1131weight : float ( 5 downto -14 ) := to_float (0.750079,5,14);

Signal ProductNode_Float1131Output_1455: float (5 downto -14);
Signal ProductNode_Float1132weight : float ( 5 downto -14 ) := to_float (0.947231,5,14);

Signal ProductNode_Float1132Output_1456: float (5 downto -14);
Signal SumNode_Float324Output_1457: float (5 downto -14);
Signal ProductNode_Float1133Output_1458: float (5 downto -14);
Signal ProductNode_Float1134weight : float ( 5 downto -14 ) := to_float (0.807766,5,14);

Signal ProductNode_Float1134Output_1459: float (5 downto -14);
Signal ProductNode_Float1135weight : float ( 5 downto -14 ) := to_float (0.825885,5,14);

Signal ProductNode_Float1135Output_1460: float (5 downto -14);
Signal ProductNode_Float1136weight : float ( 5 downto -14 ) := to_float (0.617466,5,14);

Signal ProductNode_Float1136Output_1461: float (5 downto -14);
Signal ProductNode_Float1137weight : float ( 5 downto -14 ) := to_float (0.981367,5,14);

Signal ProductNode_Float1137Output_1462: float (5 downto -14);
Signal SumNode_Float325Output_1463: float (5 downto -14);
Signal ProductNode_Float1138Output_1464: float (5 downto -14);
Signal ProductNode_Float1139weight : float ( 5 downto -14 ) := to_float (0.919167,5,14);

Signal ProductNode_Float1139Output_1465: float (5 downto -14);
Signal ProductNode_Float1140weight : float ( 5 downto -14 ) := to_float (0.933580,5,14);

Signal ProductNode_Float1140Output_1466: float (5 downto -14);
Signal SumNode_Float326Output_1467: float (5 downto -14);
Signal ProductNode_Float1141Output_1468: float (5 downto -14);
Signal SumNode_Float327Output_1469: float (5 downto -14);
Signal ProductNode_Float1142Output_1470: float (5 downto -14);
Signal ProductNode_Float1143weight : float ( 5 downto -14 ) := to_float (0.815442,5,14);

Signal ProductNode_Float1143Output_1471: float (5 downto -14);
Signal SumNode_Float328Output_1472: float (5 downto -14);
Signal ProductNode_Float1144Output_1473: float (5 downto -14);
Signal SumNode_Float329Output_1474: float (5 downto -14);
Signal ProductNode_Float1145Output_1475: float (5 downto -14);
Signal SumNode_Float330Output_1476: float (5 downto -14);
Signal ProductNode_Float1146Output_1477: float (5 downto -14);
Signal ProductNode_Float1147weight : float ( 5 downto -14 ) := to_float (0.848299,5,14);

Signal ProductNode_Float1147Output_1478: float (5 downto -14);
Signal ProductNode_Float1148weight : float ( 5 downto -14 ) := to_float (0.895308,5,14);

Signal ProductNode_Float1148Output_1479: float (5 downto -14);
Signal ProductNode_Float1149weight : float ( 5 downto -14 ) := to_float (0.842608,5,14);

Signal ProductNode_Float1149Output_1480: float (5 downto -14);
Signal SumNode_Float331Output_1481: float (5 downto -14);
Signal ProductNode_Float1150Output_1482: float (5 downto -14);
Signal ProductNode_Float1151weight : float ( 5 downto -14 ) := to_float (0.870697,5,14);

Signal ProductNode_Float1151Output_1483: float (5 downto -14);
Signal ProductNode_Float1152weight : float ( 5 downto -14 ) := to_float (0.945793,5,14);

Signal ProductNode_Float1152Output_1484: float (5 downto -14);
Signal ProductNode_Float1153weight : float ( 5 downto -14 ) := to_float (0.954870,5,14);

Signal ProductNode_Float1153Output_1485: float (5 downto -14);
Signal ProductNode_Float1154weight : float ( 5 downto -14 ) := to_float (0.870404,5,14);

Signal ProductNode_Float1154Output_1486: float (5 downto -14);
Signal ProductNode_Float1155weight : float ( 5 downto -14 ) := to_float (0.780732,5,14);

Signal ProductNode_Float1155Output_1487: float (5 downto -14);
Signal ProductNode_Float1156weight : float ( 5 downto -14 ) := to_float (0.810846,5,14);

Signal ProductNode_Float1156Output_1488: float (5 downto -14);
Signal SumNode_Float332Output_1489: float (5 downto -14);
Signal ProductNode_Float1157Output_1490: float (5 downto -14);
Signal ProductNode_Float1158weight : float ( 5 downto -14 ) := to_float (0.991361,5,14);

Signal ProductNode_Float1158Output_1491: float (5 downto -14);
Signal ProductNode_Float1159weight : float ( 5 downto -14 ) := to_float (0.669241,5,14);

Signal ProductNode_Float1159Output_1492: float (5 downto -14);
Signal ProductNode_Float1160weight : float ( 5 downto -14 ) := to_float (0.971580,5,14);

Signal ProductNode_Float1160Output_1493: float (5 downto -14);
Signal SumNode_Float333Output_1494: float (5 downto -14);
Signal ProductNode_Float1161Output_1495: float (5 downto -14);
Signal ProductNode_Float1162weight : float ( 5 downto -14 ) := to_float (0.870697,5,14);

Signal ProductNode_Float1162Output_1496: float (5 downto -14);
Signal ProductNode_Float1163weight : float ( 5 downto -14 ) := to_float (0.753690,5,14);

Signal ProductNode_Float1163Output_1497: float (5 downto -14);
Signal ProductNode_Float1164weight : float ( 5 downto -14 ) := to_float (0.774480,5,14);

Signal ProductNode_Float1164Output_1498: float (5 downto -14);
Signal ProductNode_Float1165weight : float ( 5 downto -14 ) := to_float (0.870404,5,14);

Signal ProductNode_Float1165Output_1499: float (5 downto -14);
Signal ProductNode_Float1166weight : float ( 5 downto -14 ) := to_float (0.933776,5,14);

Signal ProductNode_Float1166Output_1500: float (5 downto -14);
Signal ProductNode_Float1167weight : float ( 5 downto -14 ) := to_float (0.660973,5,14);

Signal ProductNode_Float1167Output_1501: float (5 downto -14);
Signal SumNode_Float334Output_1502: float (5 downto -14);
Signal ProductNode_Float1168Output_1503: float (5 downto -14);
Signal ProductNode_Float1169weight : float ( 5 downto -14 ) := to_float (0.870239,5,14);

Signal ProductNode_Float1169Output_1504: float (5 downto -14);
Signal SumNode_Float335Output_1505: float (5 downto -14);
Signal ProductNode_Float1170Output_1506: float (5 downto -14);
Signal ProductNode_Float1171weight : float ( 5 downto -14 ) := to_float (0.944720,5,14);

Signal ProductNode_Float1171Output_1507: float (5 downto -14);
Signal ProductNode_Float1172weight : float ( 5 downto -14 ) := to_float (0.890735,5,14);

Signal ProductNode_Float1172Output_1508: float (5 downto -14);
Signal ProductNode_Float1173weight : float ( 5 downto -14 ) := to_float (0.689002,5,14);

Signal ProductNode_Float1173Output_1509: float (5 downto -14);
Signal ProductNode_Float1174weight : float ( 5 downto -14 ) := to_float (0.966814,5,14);

Signal ProductNode_Float1174Output_1510: float (5 downto -14);
Signal SumNode_Float336Output_1511: float (5 downto -14);
Signal ProductNode_Float1175Output_1512: float (5 downto -14);
Signal ProductNode_Float1176weight : float ( 5 downto -14 ) := to_float (0.551341,5,14);

Signal ProductNode_Float1176Output_1513: float (5 downto -14);
Signal ProductNode_Float1177weight : float ( 5 downto -14 ) := to_float (0.795357,5,14);

Signal ProductNode_Float1177Output_1514: float (5 downto -14);
Signal ProductNode_Float1178weight : float ( 5 downto -14 ) := to_float (0.746308,5,14);

Signal ProductNode_Float1178Output_1515: float (5 downto -14);
Signal ProductNode_Float1179weight : float ( 5 downto -14 ) := to_float (0.989597,5,14);

Signal ProductNode_Float1179Output_1516: float (5 downto -14);
Signal ProductNode_Float1180weight : float ( 5 downto -14 ) := to_float (0.577708,5,14);

Signal ProductNode_Float1180Output_1517: float (5 downto -14);
Signal ProductNode_Float1181weight : float ( 5 downto -14 ) := to_float (0.618274,5,14);

Signal ProductNode_Float1181Output_1518: float (5 downto -14);
Signal SumNode_Float337Output_1519: float (5 downto -14);
Signal ProductNode_Float1182Output_1520: float (5 downto -14);
Signal ProductNode_Float1183weight : float ( 5 downto -14 ) := to_float (0.952809,5,14);

Signal ProductNode_Float1183Output_1521: float (5 downto -14);
Signal ProductNode_Float1184weight : float ( 5 downto -14 ) := to_float (0.495915,5,14);

Signal ProductNode_Float1184Output_1522: float (5 downto -14);
Signal ProductNode_Float1185weight : float ( 5 downto -14 ) := to_float (0.993928,5,14);

Signal ProductNode_Float1185Output_1523: float (5 downto -14);
Signal SumNode_Float338Output_1524: float (5 downto -14);
Signal ProductNode_Float1186Output_1525: float (5 downto -14);
Signal ProductNode_Float1187weight : float ( 5 downto -14 ) := to_float (0.551341,5,14);

Signal ProductNode_Float1187Output_1526: float (5 downto -14);
Signal ProductNode_Float1188weight : float ( 5 downto -14 ) := to_float (0.926235,5,14);

Signal ProductNode_Float1188Output_1527: float (5 downto -14);
Signal ProductNode_Float1189weight : float ( 5 downto -14 ) := to_float (0.616494,5,14);

Signal ProductNode_Float1189Output_1528: float (5 downto -14);
Signal ProductNode_Float1190weight : float ( 5 downto -14 ) := to_float (0.989597,5,14);

Signal ProductNode_Float1190Output_1529: float (5 downto -14);
Signal ProductNode_Float1191weight : float ( 5 downto -14 ) := to_float (0.986786,5,14);

Signal ProductNode_Float1191Output_1530: float (5 downto -14);
Signal ProductNode_Float1192weight : float ( 5 downto -14 ) := to_float (0.464416,5,14);

Signal ProductNode_Float1192Output_1531: float (5 downto -14);
Signal SumNode_Float339Output_1532: float (5 downto -14);
Signal ProductNode_Float1193Output_1533: float (5 downto -14);
Signal ProductNode_Float1194weight : float ( 5 downto -14 ) := to_float (0.770987,5,14);

Signal ProductNode_Float1194Output_1534: float (5 downto -14);
Signal SumNode_Float340Output_1535: float (5 downto -14);
Signal ProductNode_Float1195Output_1536: float (5 downto -14);
Signal ProductNode_Float1196weight : float ( 5 downto -14 ) := to_float (0.827729,5,14);

Signal ProductNode_Float1196Output_1537: float (5 downto -14);
Signal SumNode_Float341Output_1538: float (5 downto -14);
Signal ProductNode_Float1197Output_1539: float (5 downto -14);
Signal ProductNode_Float1198weight : float ( 5 downto -14 ) := to_float (0.579175,5,14);

Signal ProductNode_Float1198Output_1540: float (5 downto -14);
Signal ProductNode_Float1199weight : float ( 5 downto -14 ) := to_float (0.848299,5,14);

Signal ProductNode_Float1199Output_1541: float (5 downto -14);
Signal ProductNode_Float1200weight : float ( 5 downto -14 ) := to_float (0.562709,5,14);

Signal ProductNode_Float1200Output_1542: float (5 downto -14);
Signal ProductNode_Float1201weight : float ( 5 downto -14 ) := to_float (0.988453,5,14);

Signal ProductNode_Float1201Output_1543: float (5 downto -14);
Signal SumNode_Float342Output_1544: float (5 downto -14);
Signal ProductNode_Float1202Output_1545: float (5 downto -14);
Signal ProductNode_Float1203weight : float ( 5 downto -14 ) := to_float (0.870697,5,14);

Signal ProductNode_Float1203Output_1546: float (5 downto -14);
Signal ProductNode_Float1204weight : float ( 5 downto -14 ) := to_float (0.945793,5,14);

Signal ProductNode_Float1204Output_1547: float (5 downto -14);
Signal ProductNode_Float1205weight : float ( 5 downto -14 ) := to_float (0.729204,5,14);

Signal ProductNode_Float1205Output_1548: float (5 downto -14);
Signal ProductNode_Float1206weight : float ( 5 downto -14 ) := to_float (0.870404,5,14);

Signal ProductNode_Float1206Output_1549: float (5 downto -14);
Signal ProductNode_Float1207weight : float ( 5 downto -14 ) := to_float (0.780732,5,14);

Signal ProductNode_Float1207Output_1550: float (5 downto -14);
Signal ProductNode_Float1208weight : float ( 5 downto -14 ) := to_float (0.917308,5,14);

Signal ProductNode_Float1208Output_1551: float (5 downto -14);
Signal SumNode_Float343Output_1552: float (5 downto -14);
Signal ProductNode_Float1209Output_1553: float (5 downto -14);
Signal ProductNode_Float1210weight : float ( 5 downto -14 ) := to_float (0.979033,5,14);

Signal ProductNode_Float1210Output_1554: float (5 downto -14);
Signal ProductNode_Float1211weight : float ( 5 downto -14 ) := to_float (0.453222,5,14);

Signal ProductNode_Float1211Output_1555: float (5 downto -14);
Signal ProductNode_Float1212weight : float ( 5 downto -14 ) := to_float (0.996146,5,14);

Signal ProductNode_Float1212Output_1556: float (5 downto -14);
Signal SumNode_Float344Output_1557: float (5 downto -14);
Signal ProductNode_Float1213Output_1558: float (5 downto -14);
Signal ProductNode_Float1214weight : float ( 5 downto -14 ) := to_float (0.870697,5,14);

Signal ProductNode_Float1214Output_1559: float (5 downto -14);
Signal ProductNode_Float1215weight : float ( 5 downto -14 ) := to_float (0.753690,5,14);

Signal ProductNode_Float1215Output_1560: float (5 downto -14);
Signal ProductNode_Float1216weight : float ( 5 downto -14 ) := to_float (0.936763,5,14);

Signal ProductNode_Float1216Output_1561: float (5 downto -14);
Signal ProductNode_Float1217weight : float ( 5 downto -14 ) := to_float (0.870404,5,14);

Signal ProductNode_Float1217Output_1562: float (5 downto -14);
Signal ProductNode_Float1218weight : float ( 5 downto -14 ) := to_float (0.933776,5,14);

Signal ProductNode_Float1218Output_1563: float (5 downto -14);
Signal ProductNode_Float1219weight : float ( 5 downto -14 ) := to_float (0.973389,5,14);

Signal ProductNode_Float1219Output_1564: float (5 downto -14);
Signal SumNode_Float345Output_1565: float (5 downto -14);
Signal ProductNode_Float1220Output_1566: float (5 downto -14);
Signal ProductNode_Float1221weight : float ( 5 downto -14 ) := to_float (0.818419,5,14);

Signal ProductNode_Float1221Output_1567: float (5 downto -14);
Signal SumNode_Float346Output_1568: float (5 downto -14);
Signal ProductNode_Float1222Output_1569: float (5 downto -14);
Signal ProductNode_Float1223weight : float ( 5 downto -14 ) := to_float (0.766253,5,14);

Signal ProductNode_Float1223Output_1570: float (5 downto -14);
Signal ProductNode_Float1224weight : float ( 5 downto -14 ) := to_float (0.890735,5,14);

Signal ProductNode_Float1224Output_1571: float (5 downto -14);
Signal ProductNode_Float1225weight : float ( 5 downto -14 ) := to_float (0.382644,5,14);

Signal ProductNode_Float1225Output_1572: float (5 downto -14);
Signal ProductNode_Float1226weight : float ( 5 downto -14 ) := to_float (0.998354,5,14);

Signal ProductNode_Float1226Output_1573: float (5 downto -14);
Signal SumNode_Float347Output_1574: float (5 downto -14);
Signal ProductNode_Float1227Output_1575: float (5 downto -14);
Signal ProductNode_Float1228weight : float ( 5 downto -14 ) := to_float (0.551341,5,14);

Signal ProductNode_Float1228Output_1576: float (5 downto -14);
Signal ProductNode_Float1229weight : float ( 5 downto -14 ) := to_float (0.795357,5,14);

Signal ProductNode_Float1229Output_1577: float (5 downto -14);
Signal ProductNode_Float1230weight : float ( 5 downto -14 ) := to_float (0.948695,5,14);

Signal ProductNode_Float1230Output_1578: float (5 downto -14);
Signal ProductNode_Float1231weight : float ( 5 downto -14 ) := to_float (0.989597,5,14);

Signal ProductNode_Float1231Output_1579: float (5 downto -14);
Signal ProductNode_Float1232weight : float ( 5 downto -14 ) := to_float (0.577708,5,14);

Signal ProductNode_Float1232Output_1580: float (5 downto -14);
Signal ProductNode_Float1233weight : float ( 5 downto -14 ) := to_float (0.981240,5,14);

Signal ProductNode_Float1233Output_1581: float (5 downto -14);
Signal SumNode_Float348Output_1582: float (5 downto -14);
Signal ProductNode_Float1234Output_1583: float (5 downto -14);
Signal ProductNode_Float1235weight : float ( 5 downto -14 ) := to_float (0.960334,5,14);

Signal ProductNode_Float1235Output_1584: float (5 downto -14);
Signal ProductNode_Float1236weight : float ( 5 downto -14 ) := to_float (0.336149,5,14);

Signal ProductNode_Float1236Output_1585: float (5 downto -14);
Signal ProductNode_Float1237weight : float ( 5 downto -14 ) := to_float (0.999140,5,14);

Signal ProductNode_Float1237Output_1586: float (5 downto -14);
Signal SumNode_Float349Output_1587: float (5 downto -14);
Signal ProductNode_Float1238Output_1588: float (5 downto -14);
Signal ProductNode_Float1239weight : float ( 5 downto -14 ) := to_float (0.551341,5,14);

Signal ProductNode_Float1239Output_1589: float (5 downto -14);
Signal ProductNode_Float1240weight : float ( 5 downto -14 ) := to_float (0.926235,5,14);

Signal ProductNode_Float1240Output_1590: float (5 downto -14);
Signal ProductNode_Float1241weight : float ( 5 downto -14 ) := to_float (0.981519,5,14);

Signal ProductNode_Float1241Output_1591: float (5 downto -14);
Signal ProductNode_Float1242weight : float ( 5 downto -14 ) := to_float (0.989597,5,14);

Signal ProductNode_Float1242Output_1592: float (5 downto -14);
Signal ProductNode_Float1243weight : float ( 5 downto -14 ) := to_float (0.986786,5,14);

Signal ProductNode_Float1243Output_1593: float (5 downto -14);
Signal ProductNode_Float1244weight : float ( 5 downto -14 ) := to_float (0.995641,5,14);

Signal ProductNode_Float1244Output_1594: float (5 downto -14);
Signal SumNode_Float350Output_1595: float (5 downto -14);
Signal ProductNode_Float1245Output_1596: float (5 downto -14);
Signal ProductNode_Float1246weight : float ( 5 downto -14 ) := to_float (0.664315,5,14);

Signal ProductNode_Float1246Output_1597: float (5 downto -14);
Signal SumNode_Float351Output_1598: float (5 downto -14);
Signal ProductNode_Float1247Output_1599: float (5 downto -14);
Signal ProductNode_Float1248weight : float ( 5 downto -14 ) := to_float (0.634118,5,14);

Signal ProductNode_Float1248Output_1600: float (5 downto -14);
Signal SumNode_Float352Output_1601: float (5 downto -14);
Signal ProductNode_Float1249Output_1602: float (5 downto -14);
Signal ProductNode_Float1250weight : float ( 5 downto -14 ) := to_float (0.760169,5,14);

Signal ProductNode_Float1250Output_1603: float (5 downto -14);
Signal SumNode_Float353Output_1604: float (5 downto -14);
Signal ProductNode_Float1251Output_1605: float (5 downto -14);
Signal ProductNode_Float1252weight : float ( 5 downto -14 ) := to_float (0.970921,5,14);

Signal ProductNode_Float1252Output_1606: float (5 downto -14);
Signal ProductNode_Float1253weight : float ( 5 downto -14 ) := to_float (0.672140,5,14);

Signal ProductNode_Float1253Output_1607: float (5 downto -14);
Signal SumNode_Float354Output_1608: float (5 downto -14);
Signal ProductNode_Float1254Output_1609: float (5 downto -14);
Signal ProductNode_Float1255weight : float ( 5 downto -14 ) := to_float (0.989270,5,14);

Signal ProductNode_Float1255Output_1610: float (5 downto -14);
Signal ProductNode_Float1256weight : float ( 5 downto -14 ) := to_float (0.997554,5,14);

Signal ProductNode_Float1256Output_1611: float (5 downto -14);
Signal ProductNode_Float1257weight : float ( 5 downto -14 ) := to_float (0.414069,5,14);

Signal ProductNode_Float1257Output_1612: float (5 downto -14);
Signal SumNode_Float355Output_1613: float (5 downto -14);
Signal ProductNode_Float1258Output_1614: float (5 downto -14);
Signal ProductNode_Float1259weight : float ( 5 downto -14 ) := to_float (0.853307,5,14);

Signal ProductNode_Float1259Output_1615: float (5 downto -14);
Signal ProductNode_Float1260weight : float ( 5 downto -14 ) := to_float (0.886527,5,14);

Signal ProductNode_Float1260Output_1616: float (5 downto -14);
Signal SumNode_Float356Output_1617: float (5 downto -14);
Signal ProductNode_Float1261Output_1618: float (5 downto -14);
Signal ProductNode_Float1262weight : float ( 5 downto -14 ) := to_float (0.554692,5,14);

Signal ProductNode_Float1262Output_1619: float (5 downto -14);
Signal ProductNode_Float1263weight : float ( 5 downto -14 ) := to_float (0.989739,5,14);

Signal ProductNode_Float1263Output_1620: float (5 downto -14);
Signal ProductNode_Float1264weight : float ( 5 downto -14 ) := to_float (0.549861,5,14);

Signal ProductNode_Float1264Output_1621: float (5 downto -14);
Signal SumNode_Float357Output_1622: float (5 downto -14);
Signal ProductNode_Float1265Output_1623: float (5 downto -14);
Signal SumNode_Float358Output_1624: float (5 downto -14);
Signal ProductNode_Float1266Output_1625: float (5 downto -14);
Signal ProductNode_Float1267weight : float ( 5 downto -14 ) := to_float (0.994862,5,14);

Signal ProductNode_Float1267Output_1626: float (5 downto -14);
Signal ProductNode_Float1268weight : float ( 5 downto -14 ) := to_float (0.817897,5,14);

Signal ProductNode_Float1268Output_1627: float (5 downto -14);
Signal ProductNode_Float1269weight : float ( 5 downto -14 ) := to_float (0.912886,5,14);

Signal ProductNode_Float1269Output_1628: float (5 downto -14);
Signal SumNode_Float359Output_1629: float (5 downto -14);
Signal ProductNode_Float1270Output_1630: float (5 downto -14);
Signal ProductNode_Float1271weight : float ( 5 downto -14 ) := to_float (0.976301,5,14);

Signal ProductNode_Float1271Output_1631: float (5 downto -14);
Signal ProductNode_Float1272weight : float ( 5 downto -14 ) := to_float (0.988880,5,14);

Signal ProductNode_Float1272Output_1632: float (5 downto -14);
Signal ProductNode_Float1273weight : float ( 5 downto -14 ) := to_float (0.558577,5,14);

Signal ProductNode_Float1273Output_1633: float (5 downto -14);
Signal SumNode_Float360Output_1634: float (5 downto -14);
Signal ProductNode_Float1274Output_1635: float (5 downto -14);
Signal ProductNode_Float1275weight : float ( 5 downto -14 ) := to_float (0.731617,5,14);

Signal ProductNode_Float1275Output_1636: float (5 downto -14);
Signal ProductNode_Float1276weight : float ( 5 downto -14 ) := to_float (0.954043,5,14);

Signal ProductNode_Float1276Output_1637: float (5 downto -14);
Signal SumNode_Float361Output_1638: float (5 downto -14);
Signal ProductNode_Float1277Output_1639: float (5 downto -14);
Signal ProductNode_Float1278weight : float ( 5 downto -14 ) := to_float (0.646579,5,14);

Signal ProductNode_Float1278Output_1640: float (5 downto -14);
Signal ProductNode_Float1279weight : float ( 5 downto -14 ) := to_float (0.985013,5,14);

Signal ProductNode_Float1279Output_1641: float (5 downto -14);
Signal ProductNode_Float1280weight : float ( 5 downto -14 ) := to_float (0.592017,5,14);

Signal ProductNode_Float1280Output_1642: float (5 downto -14);
Signal SumNode_Float362Output_1643: float (5 downto -14);
Signal ProductNode_Float1281Output_1644: float (5 downto -14);
Signal SumNode_Float363Output_1645: float (5 downto -14);
Signal ProductNode_Float1282Output_1646: float (5 downto -14);
Signal ProductNode_Float1283weight : float ( 5 downto -14 ) := to_float (0.479802,5,14);

Signal ProductNode_Float1283Output_1647: float (5 downto -14);
Signal SumNode_Float364Output_1648: float (5 downto -14);
Signal ProductNode_Float1284Output_1649: float (5 downto -14);
Signal ProductNode_Float1285weight : float ( 5 downto -14 ) := to_float (0.807423,5,14);

Signal ProductNode_Float1285Output_1650: float (5 downto -14);
Signal ProductNode_Float1286weight : float ( 5 downto -14 ) := to_float (0.919372,5,14);

Signal ProductNode_Float1286Output_1651: float (5 downto -14);
Signal SumNode_Float365Output_1652: float (5 downto -14);
Signal ProductNode_Float1287Output_1653: float (5 downto -14);
Signal ProductNode_Float1288weight : float ( 5 downto -14 ) := to_float (0.694473,5,14);

Signal ProductNode_Float1288Output_1654: float (5 downto -14);
Signal ProductNode_Float1289weight : float ( 5 downto -14 ) := to_float (0.843444,5,14);

Signal ProductNode_Float1289Output_1655: float (5 downto -14);
Signal ProductNode_Float1290weight : float ( 5 downto -14 ) := to_float (0.682797,5,14);

Signal ProductNode_Float1290Output_1656: float (5 downto -14);
Signal ProductNode_Float1291weight : float ( 5 downto -14 ) := to_float (0.968381,5,14);

Signal ProductNode_Float1291Output_1657: float (5 downto -14);
Signal SumNode_Float366Output_1658: float (5 downto -14);
Signal ProductNode_Float1292Output_1659: float (5 downto -14);
Signal ProductNode_Float1293weight : float ( 5 downto -14 ) := to_float (0.965376,5,14);

Signal ProductNode_Float1293Output_1660: float (5 downto -14);
Signal ProductNode_Float1294weight : float ( 5 downto -14 ) := to_float (0.697447,5,14);

Signal ProductNode_Float1294Output_1661: float (5 downto -14);
Signal SumNode_Float367Output_1662: float (5 downto -14);
Signal ProductNode_Float1295Output_1663: float (5 downto -14);
Signal ProductNode_Float1296weight : float ( 5 downto -14 ) := to_float (0.970921,5,14);

Signal ProductNode_Float1296Output_1664: float (5 downto -14);
Signal ProductNode_Float1297weight : float ( 5 downto -14 ) := to_float (0.672140,5,14);

Signal ProductNode_Float1297Output_1665: float (5 downto -14);
Signal SumNode_Float368Output_1666: float (5 downto -14);
Signal ProductNode_Float1298Output_1667: float (5 downto -14);
Signal ProductNode_Float1299weight : float ( 5 downto -14 ) := to_float (0.989270,5,14);

Signal ProductNode_Float1299Output_1668: float (5 downto -14);
Signal ProductNode_Float1300weight : float ( 5 downto -14 ) := to_float (0.997554,5,14);

Signal ProductNode_Float1300Output_1669: float (5 downto -14);
Signal ProductNode_Float1301weight : float ( 5 downto -14 ) := to_float (0.414069,5,14);

Signal ProductNode_Float1301Output_1670: float (5 downto -14);
Signal SumNode_Float369Output_1671: float (5 downto -14);
Signal ProductNode_Float1302Output_1672: float (5 downto -14);
Signal ProductNode_Float1303weight : float ( 5 downto -14 ) := to_float (0.853307,5,14);

Signal ProductNode_Float1303Output_1673: float (5 downto -14);
Signal ProductNode_Float1304weight : float ( 5 downto -14 ) := to_float (0.886527,5,14);

Signal ProductNode_Float1304Output_1674: float (5 downto -14);
Signal SumNode_Float370Output_1675: float (5 downto -14);
Signal ProductNode_Float1305Output_1676: float (5 downto -14);
Signal ProductNode_Float1306weight : float ( 5 downto -14 ) := to_float (0.554692,5,14);

Signal ProductNode_Float1306Output_1677: float (5 downto -14);
Signal ProductNode_Float1307weight : float ( 5 downto -14 ) := to_float (0.989739,5,14);

Signal ProductNode_Float1307Output_1678: float (5 downto -14);
Signal ProductNode_Float1308weight : float ( 5 downto -14 ) := to_float (0.549861,5,14);

Signal ProductNode_Float1308Output_1679: float (5 downto -14);
Signal SumNode_Float371Output_1680: float (5 downto -14);
Signal ProductNode_Float1309Output_1681: float (5 downto -14);
Signal SumNode_Float372Output_1682: float (5 downto -14);
Signal ProductNode_Float1310Output_1683: float (5 downto -14);
Signal ProductNode_Float1311weight : float ( 5 downto -14 ) := to_float (0.970629,5,14);

Signal ProductNode_Float1311Output_1684: float (5 downto -14);
Signal ProductNode_Float1312weight : float ( 5 downto -14 ) := to_float (0.817897,5,14);

Signal ProductNode_Float1312Output_1685: float (5 downto -14);
Signal ProductNode_Float1313weight : float ( 5 downto -14 ) := to_float (0.912886,5,14);

Signal ProductNode_Float1313Output_1686: float (5 downto -14);
Signal SumNode_Float373Output_1687: float (5 downto -14);
Signal ProductNode_Float1314Output_1688: float (5 downto -14);
Signal ProductNode_Float1315weight : float ( 5 downto -14 ) := to_float (0.976301,5,14);

Signal ProductNode_Float1315Output_1689: float (5 downto -14);
Signal ProductNode_Float1316weight : float ( 5 downto -14 ) := to_float (0.988880,5,14);

Signal ProductNode_Float1316Output_1690: float (5 downto -14);
Signal ProductNode_Float1317weight : float ( 5 downto -14 ) := to_float (0.558577,5,14);

Signal ProductNode_Float1317Output_1691: float (5 downto -14);
Signal SumNode_Float374Output_1692: float (5 downto -14);
Signal ProductNode_Float1318Output_1693: float (5 downto -14);
Signal ProductNode_Float1319weight : float ( 5 downto -14 ) := to_float (0.731617,5,14);

Signal ProductNode_Float1319Output_1694: float (5 downto -14);
Signal ProductNode_Float1320weight : float ( 5 downto -14 ) := to_float (0.954043,5,14);

Signal ProductNode_Float1320Output_1695: float (5 downto -14);
Signal SumNode_Float375Output_1696: float (5 downto -14);
Signal ProductNode_Float1321Output_1697: float (5 downto -14);
Signal ProductNode_Float1322weight : float ( 5 downto -14 ) := to_float (0.646579,5,14);

Signal ProductNode_Float1322Output_1698: float (5 downto -14);
Signal ProductNode_Float1323weight : float ( 5 downto -14 ) := to_float (0.985013,5,14);

Signal ProductNode_Float1323Output_1699: float (5 downto -14);
Signal ProductNode_Float1324weight : float ( 5 downto -14 ) := to_float (0.592017,5,14);

Signal ProductNode_Float1324Output_1700: float (5 downto -14);
Signal SumNode_Float376Output_1701: float (5 downto -14);
Signal ProductNode_Float1325Output_1702: float (5 downto -14);
Signal SumNode_Float377Output_1703: float (5 downto -14);
Signal ProductNode_Float1326Output_1704: float (5 downto -14);
Signal ProductNode_Float1327weight : float ( 5 downto -14 ) := to_float (0.673404,5,14);

Signal ProductNode_Float1327Output_1705: float (5 downto -14);
Signal SumNode_Float378Output_1706: float (5 downto -14);
Signal ProductNode_Float1328Output_1707: float (5 downto -14);
Signal ProductNode_Float1329weight : float ( 5 downto -14 ) := to_float (0.623360,5,14);

Signal ProductNode_Float1329Output_1708: float (5 downto -14);
Signal ProductNode_Float1330weight : float ( 5 downto -14 ) := to_float (0.980424,5,14);

Signal ProductNode_Float1330Output_1709: float (5 downto -14);
Signal SumNode_Float379Output_1710: float (5 downto -14);
Signal ProductNode_Float1331Output_1711: float (5 downto -14);
Signal ProductNode_Float1332weight : float ( 5 downto -14 ) := to_float (0.694473,5,14);

Signal ProductNode_Float1332Output_1712: float (5 downto -14);
Signal ProductNode_Float1333weight : float ( 5 downto -14 ) := to_float (0.894649,5,14);

Signal ProductNode_Float1333Output_1713: float (5 downto -14);
Signal ProductNode_Float1334weight : float ( 5 downto -14 ) := to_float (0.482891,5,14);

Signal ProductNode_Float1334Output_1714: float (5 downto -14);
Signal ProductNode_Float1335weight : float ( 5 downto -14 ) := to_float (0.994693,5,14);

Signal ProductNode_Float1335Output_1715: float (5 downto -14);
Signal SumNode_Float380Output_1716: float (5 downto -14);
Signal ProductNode_Float1336Output_1717: float (5 downto -14);
Signal ProductNode_Float1337weight : float ( 5 downto -14 ) := to_float (0.965376,5,14);

Signal ProductNode_Float1337Output_1718: float (5 downto -14);
Signal ProductNode_Float1338weight : float ( 5 downto -14 ) := to_float (0.964572,5,14);

Signal ProductNode_Float1338Output_1719: float (5 downto -14);
Signal SumNode_Float381Output_1720: float (5 downto -14);
Signal ProductNode_Float1339Output_1721: float (5 downto -14);
Signal SumNode_Float382Output_1722: float (5 downto -14);
Signal ProductNode_Float1340Output_1723: float (5 downto -14);
Signal ProductNode_Float1341weight : float ( 5 downto -14 ) := to_float (0.952231,5,14);

Signal ProductNode_Float1341Output_1724: float (5 downto -14);
Signal ProductNode_Float1342weight : float ( 5 downto -14 ) := to_float (0.970921,5,14);

Signal ProductNode_Float1342Output_1725: float (5 downto -14);
Signal ProductNode_Float1343weight : float ( 5 downto -14 ) := to_float (0.672140,5,14);

Signal ProductNode_Float1343Output_1726: float (5 downto -14);
Signal SumNode_Float383Output_1727: float (5 downto -14);
Signal ProductNode_Float1344Output_1728: float (5 downto -14);
Signal ProductNode_Float1345weight : float ( 5 downto -14 ) := to_float (0.989270,5,14);

Signal ProductNode_Float1345Output_1729: float (5 downto -14);
Signal ProductNode_Float1346weight : float ( 5 downto -14 ) := to_float (0.966381,5,14);

Signal ProductNode_Float1346Output_1730: float (5 downto -14);
Signal ProductNode_Float1347weight : float ( 5 downto -14 ) := to_float (0.690672,5,14);

Signal ProductNode_Float1347Output_1731: float (5 downto -14);
Signal SumNode_Float384Output_1732: float (5 downto -14);
Signal ProductNode_Float1348Output_1733: float (5 downto -14);
Signal ProductNode_Float1349weight : float ( 5 downto -14 ) := to_float (0.853307,5,14);

Signal ProductNode_Float1349Output_1734: float (5 downto -14);
Signal ProductNode_Float1350weight : float ( 5 downto -14 ) := to_float (0.886527,5,14);

Signal ProductNode_Float1350Output_1735: float (5 downto -14);
Signal SumNode_Float385Output_1736: float (5 downto -14);
Signal ProductNode_Float1351Output_1737: float (5 downto -14);
Signal ProductNode_Float1352weight : float ( 5 downto -14 ) := to_float (0.554692,5,14);

Signal ProductNode_Float1352Output_1738: float (5 downto -14);
Signal ProductNode_Float1353weight : float ( 5 downto -14 ) := to_float (0.941870,5,14);

Signal ProductNode_Float1353Output_1739: float (5 downto -14);
Signal ProductNode_Float1354weight : float ( 5 downto -14 ) := to_float (0.763101,5,14);

Signal ProductNode_Float1354Output_1740: float (5 downto -14);
Signal SumNode_Float386Output_1741: float (5 downto -14);
Signal ProductNode_Float1355Output_1742: float (5 downto -14);
Signal SumNode_Float387Output_1743: float (5 downto -14);
Signal ProductNode_Float1356Output_1744: float (5 downto -14);
Signal ProductNode_Float1357weight : float ( 5 downto -14 ) := to_float (0.951966,5,14);

Signal ProductNode_Float1357Output_1745: float (5 downto -14);
Signal ProductNode_Float1358weight : float ( 5 downto -14 ) := to_float (0.817897,5,14);

Signal ProductNode_Float1358Output_1746: float (5 downto -14);
Signal ProductNode_Float1359weight : float ( 5 downto -14 ) := to_float (0.912886,5,14);

Signal ProductNode_Float1359Output_1747: float (5 downto -14);
Signal SumNode_Float388Output_1748: float (5 downto -14);
Signal ProductNode_Float1360Output_1749: float (5 downto -14);
Signal ProductNode_Float1361weight : float ( 5 downto -14 ) := to_float (0.976301,5,14);

Signal ProductNode_Float1361Output_1750: float (5 downto -14);
Signal ProductNode_Float1362weight : float ( 5 downto -14 ) := to_float (0.909585,5,14);

Signal ProductNode_Float1362Output_1751: float (5 downto -14);
Signal ProductNode_Float1363weight : float ( 5 downto -14 ) := to_float (0.822920,5,14);

Signal ProductNode_Float1363Output_1752: float (5 downto -14);
Signal SumNode_Float389Output_1753: float (5 downto -14);
Signal ProductNode_Float1364Output_1754: float (5 downto -14);
Signal ProductNode_Float1365weight : float ( 5 downto -14 ) := to_float (0.731617,5,14);

Signal ProductNode_Float1365Output_1755: float (5 downto -14);
Signal ProductNode_Float1366weight : float ( 5 downto -14 ) := to_float (0.954043,5,14);

Signal ProductNode_Float1366Output_1756: float (5 downto -14);
Signal SumNode_Float390Output_1757: float (5 downto -14);
Signal ProductNode_Float1367Output_1758: float (5 downto -14);
Signal ProductNode_Float1368weight : float ( 5 downto -14 ) := to_float (0.646579,5,14);

Signal ProductNode_Float1368Output_1759: float (5 downto -14);
Signal ProductNode_Float1369weight : float ( 5 downto -14 ) := to_float (0.790147,5,14);

Signal ProductNode_Float1369Output_1760: float (5 downto -14);
Signal ProductNode_Float1370weight : float ( 5 downto -14 ) := to_float (0.929014,5,14);

Signal ProductNode_Float1370Output_1761: float (5 downto -14);
Signal SumNode_Float391Output_1762: float (5 downto -14);
Signal ProductNode_Float1371Output_1763: float (5 downto -14);
Signal SumNode_Float392Output_1764: float (5 downto -14);
Signal ProductNode_Float1372Output_1765: float (5 downto -14);
Signal ProductNode_Float1373weight : float ( 5 downto -14 ) := to_float (0.737500,5,14);

Signal ProductNode_Float1373Output_1766: float (5 downto -14);
Signal SumNode_Float393Output_1767: float (5 downto -14);
Signal ProductNode_Float1374Output_1768: float (5 downto -14);
Signal ProductNode_Float1375weight : float ( 5 downto -14 ) := to_float (0.807423,5,14);

Signal ProductNode_Float1375Output_1769: float (5 downto -14);
Signal ProductNode_Float1376weight : float ( 5 downto -14 ) := to_float (0.919372,5,14);

Signal ProductNode_Float1376Output_1770: float (5 downto -14);
Signal SumNode_Float394Output_1771: float (5 downto -14);
Signal ProductNode_Float1377Output_1772: float (5 downto -14);
Signal ProductNode_Float1378weight : float ( 5 downto -14 ) := to_float (0.579487,5,14);

Signal ProductNode_Float1378Output_1773: float (5 downto -14);
Signal ProductNode_Float1379weight : float ( 5 downto -14 ) := to_float (0.790558,5,14);

Signal ProductNode_Float1379Output_1774: float (5 downto -14);
Signal ProductNode_Float1380weight : float ( 5 downto -14 ) := to_float (0.682797,5,14);

Signal ProductNode_Float1380Output_1775: float (5 downto -14);
Signal ProductNode_Float1381weight : float ( 5 downto -14 ) := to_float (0.968381,5,14);

Signal ProductNode_Float1381Output_1776: float (5 downto -14);
Signal SumNode_Float395Output_1777: float (5 downto -14);
Signal ProductNode_Float1382Output_1778: float (5 downto -14);
Signal ProductNode_Float1383weight : float ( 5 downto -14 ) := to_float (0.986575,5,14);

Signal ProductNode_Float1383Output_1779: float (5 downto -14);
Signal ProductNode_Float1384weight : float ( 5 downto -14 ) := to_float (0.578242,5,14);

Signal ProductNode_Float1384Output_1780: float (5 downto -14);
Signal SumNode_Float396Output_1781: float (5 downto -14);
Signal ProductNode_Float1385Output_1782: float (5 downto -14);
Signal ProductNode_Float1386weight : float ( 5 downto -14 ) := to_float (0.970921,5,14);

Signal ProductNode_Float1386Output_1783: float (5 downto -14);
Signal ProductNode_Float1387weight : float ( 5 downto -14 ) := to_float (0.672140,5,14);

Signal ProductNode_Float1387Output_1784: float (5 downto -14);
Signal SumNode_Float397Output_1785: float (5 downto -14);
Signal ProductNode_Float1388Output_1786: float (5 downto -14);
Signal ProductNode_Float1389weight : float ( 5 downto -14 ) := to_float (0.989270,5,14);

Signal ProductNode_Float1389Output_1787: float (5 downto -14);
Signal ProductNode_Float1390weight : float ( 5 downto -14 ) := to_float (0.966381,5,14);

Signal ProductNode_Float1390Output_1788: float (5 downto -14);
Signal ProductNode_Float1391weight : float ( 5 downto -14 ) := to_float (0.690672,5,14);

Signal ProductNode_Float1391Output_1789: float (5 downto -14);
Signal SumNode_Float398Output_1790: float (5 downto -14);
Signal ProductNode_Float1392Output_1791: float (5 downto -14);
Signal ProductNode_Float1393weight : float ( 5 downto -14 ) := to_float (0.853307,5,14);

Signal ProductNode_Float1393Output_1792: float (5 downto -14);
Signal ProductNode_Float1394weight : float ( 5 downto -14 ) := to_float (0.886527,5,14);

Signal ProductNode_Float1394Output_1793: float (5 downto -14);
Signal SumNode_Float399Output_1794: float (5 downto -14);
Signal ProductNode_Float1395Output_1795: float (5 downto -14);
Signal ProductNode_Float1396weight : float ( 5 downto -14 ) := to_float (0.554692,5,14);

Signal ProductNode_Float1396Output_1796: float (5 downto -14);
Signal ProductNode_Float1397weight : float ( 5 downto -14 ) := to_float (0.941870,5,14);

Signal ProductNode_Float1397Output_1797: float (5 downto -14);
Signal ProductNode_Float1398weight : float ( 5 downto -14 ) := to_float (0.763101,5,14);

Signal ProductNode_Float1398Output_1798: float (5 downto -14);
Signal SumNode_Float400Output_1799: float (5 downto -14);
Signal ProductNode_Float1399Output_1800: float (5 downto -14);
Signal SumNode_Float401Output_1801: float (5 downto -14);
Signal ProductNode_Float1400Output_1802: float (5 downto -14);
Signal ProductNode_Float1401weight : float ( 5 downto -14 ) := to_float (0.840616,5,14);

Signal ProductNode_Float1401Output_1803: float (5 downto -14);
Signal ProductNode_Float1402weight : float ( 5 downto -14 ) := to_float (0.817897,5,14);

Signal ProductNode_Float1402Output_1804: float (5 downto -14);
Signal ProductNode_Float1403weight : float ( 5 downto -14 ) := to_float (0.912886,5,14);

Signal ProductNode_Float1403Output_1805: float (5 downto -14);
Signal SumNode_Float402Output_1806: float (5 downto -14);
Signal ProductNode_Float1404Output_1807: float (5 downto -14);
Signal ProductNode_Float1405weight : float ( 5 downto -14 ) := to_float (0.976301,5,14);

Signal ProductNode_Float1405Output_1808: float (5 downto -14);
Signal ProductNode_Float1406weight : float ( 5 downto -14 ) := to_float (0.909585,5,14);

Signal ProductNode_Float1406Output_1809: float (5 downto -14);
Signal ProductNode_Float1407weight : float ( 5 downto -14 ) := to_float (0.822920,5,14);

Signal ProductNode_Float1407Output_1810: float (5 downto -14);
Signal SumNode_Float403Output_1811: float (5 downto -14);
Signal ProductNode_Float1408Output_1812: float (5 downto -14);
Signal ProductNode_Float1409weight : float ( 5 downto -14 ) := to_float (0.731617,5,14);

Signal ProductNode_Float1409Output_1813: float (5 downto -14);
Signal ProductNode_Float1410weight : float ( 5 downto -14 ) := to_float (0.954043,5,14);

Signal ProductNode_Float1410Output_1814: float (5 downto -14);
Signal SumNode_Float404Output_1815: float (5 downto -14);
Signal ProductNode_Float1411Output_1816: float (5 downto -14);
Signal ProductNode_Float1412weight : float ( 5 downto -14 ) := to_float (0.646579,5,14);

Signal ProductNode_Float1412Output_1817: float (5 downto -14);
Signal ProductNode_Float1413weight : float ( 5 downto -14 ) := to_float (0.790147,5,14);

Signal ProductNode_Float1413Output_1818: float (5 downto -14);
Signal ProductNode_Float1414weight : float ( 5 downto -14 ) := to_float (0.929014,5,14);

Signal ProductNode_Float1414Output_1819: float (5 downto -14);
Signal SumNode_Float405Output_1820: float (5 downto -14);
Signal ProductNode_Float1415Output_1821: float (5 downto -14);
Signal SumNode_Float406Output_1822: float (5 downto -14);
Signal ProductNode_Float1416Output_1823: float (5 downto -14);
Signal ProductNode_Float1417weight : float ( 5 downto -14 ) := to_float (0.896858,5,14);

Signal ProductNode_Float1417Output_1824: float (5 downto -14);
Signal SumNode_Float407Output_1825: float (5 downto -14);
Signal ProductNode_Float1418Output_1826: float (5 downto -14);
Signal ProductNode_Float1419weight : float ( 5 downto -14 ) := to_float (0.623360,5,14);

Signal ProductNode_Float1419Output_1827: float (5 downto -14);
Signal ProductNode_Float1420weight : float ( 5 downto -14 ) := to_float (0.980424,5,14);

Signal ProductNode_Float1420Output_1828: float (5 downto -14);
Signal SumNode_Float408Output_1829: float (5 downto -14);
Signal ProductNode_Float1421Output_1830: float (5 downto -14);
Signal ProductNode_Float1422weight : float ( 5 downto -14 ) := to_float (0.579487,5,14);

Signal ProductNode_Float1422Output_1831: float (5 downto -14);
Signal ProductNode_Float1423weight : float ( 5 downto -14 ) := to_float (0.928799,5,14);

Signal ProductNode_Float1423Output_1832: float (5 downto -14);
Signal ProductNode_Float1424weight : float ( 5 downto -14 ) := to_float (0.482891,5,14);

Signal ProductNode_Float1424Output_1833: float (5 downto -14);
Signal ProductNode_Float1425weight : float ( 5 downto -14 ) := to_float (0.994693,5,14);

Signal ProductNode_Float1425Output_1834: float (5 downto -14);
Signal SumNode_Float409Output_1835: float (5 downto -14);
Signal ProductNode_Float1426Output_1836: float (5 downto -14);
Signal ProductNode_Float1427weight : float ( 5 downto -14 ) := to_float (0.986575,5,14);

Signal ProductNode_Float1427Output_1837: float (5 downto -14);
Signal ProductNode_Float1428weight : float ( 5 downto -14 ) := to_float (0.986723,5,14);

Signal ProductNode_Float1428Output_1838: float (5 downto -14);
Signal SumNode_Float410Output_1839: float (5 downto -14);
Signal ProductNode_Float1429Output_1840: float (5 downto -14);
Signal SumNode_Float411Output_1841: float (5 downto -14);
Signal ProductNode_Float1430Output_1842: float (5 downto -14);
Signal ProductNode_Float1431weight : float ( 5 downto -14 ) := to_float (0.736765,5,14);

Signal ProductNode_Float1431Output_1843: float (5 downto -14);
Signal SumNode_Float412Output_1844: float (5 downto -14);
Signal ProductNode_Float1432Output_1845: float (5 downto -14);
Signal ProductNode_Float1433weight : float ( 5 downto -14 ) := to_float (0.848299,5,14);

Signal ProductNode_Float1433Output_1846: float (5 downto -14);
Signal ProductNode_Float1434weight : float ( 5 downto -14 ) := to_float (0.895308,5,14);

Signal ProductNode_Float1434Output_1847: float (5 downto -14);
Signal ProductNode_Float1435weight : float ( 5 downto -14 ) := to_float (0.842608,5,14);

Signal ProductNode_Float1435Output_1848: float (5 downto -14);
Signal SumNode_Float413Output_1849: float (5 downto -14);
Signal ProductNode_Float1436Output_1850: float (5 downto -14);
Signal ProductNode_Float1437weight : float ( 5 downto -14 ) := to_float (0.870697,5,14);

Signal ProductNode_Float1437Output_1851: float (5 downto -14);
Signal ProductNode_Float1438weight : float ( 5 downto -14 ) := to_float (0.945793,5,14);

Signal ProductNode_Float1438Output_1852: float (5 downto -14);
Signal ProductNode_Float1439weight : float ( 5 downto -14 ) := to_float (0.954870,5,14);

Signal ProductNode_Float1439Output_1853: float (5 downto -14);
Signal ProductNode_Float1440weight : float ( 5 downto -14 ) := to_float (0.870404,5,14);

Signal ProductNode_Float1440Output_1854: float (5 downto -14);
Signal ProductNode_Float1441weight : float ( 5 downto -14 ) := to_float (0.780732,5,14);

Signal ProductNode_Float1441Output_1855: float (5 downto -14);
Signal ProductNode_Float1442weight : float ( 5 downto -14 ) := to_float (0.810846,5,14);

Signal ProductNode_Float1442Output_1856: float (5 downto -14);
Signal SumNode_Float414Output_1857: float (5 downto -14);
Signal ProductNode_Float1443Output_1858: float (5 downto -14);
Signal ProductNode_Float1444weight : float ( 5 downto -14 ) := to_float (0.991361,5,14);

Signal ProductNode_Float1444Output_1859: float (5 downto -14);
Signal ProductNode_Float1445weight : float ( 5 downto -14 ) := to_float (0.669241,5,14);

Signal ProductNode_Float1445Output_1860: float (5 downto -14);
Signal ProductNode_Float1446weight : float ( 5 downto -14 ) := to_float (0.971580,5,14);

Signal ProductNode_Float1446Output_1861: float (5 downto -14);
Signal SumNode_Float415Output_1862: float (5 downto -14);
Signal ProductNode_Float1447Output_1863: float (5 downto -14);
Signal ProductNode_Float1448weight : float ( 5 downto -14 ) := to_float (0.870697,5,14);

Signal ProductNode_Float1448Output_1864: float (5 downto -14);
Signal ProductNode_Float1449weight : float ( 5 downto -14 ) := to_float (0.753690,5,14);

Signal ProductNode_Float1449Output_1865: float (5 downto -14);
Signal ProductNode_Float1450weight : float ( 5 downto -14 ) := to_float (0.774480,5,14);

Signal ProductNode_Float1450Output_1866: float (5 downto -14);
Signal ProductNode_Float1451weight : float ( 5 downto -14 ) := to_float (0.870404,5,14);

Signal ProductNode_Float1451Output_1867: float (5 downto -14);
Signal ProductNode_Float1452weight : float ( 5 downto -14 ) := to_float (0.933776,5,14);

Signal ProductNode_Float1452Output_1868: float (5 downto -14);
Signal ProductNode_Float1453weight : float ( 5 downto -14 ) := to_float (0.660973,5,14);

Signal ProductNode_Float1453Output_1869: float (5 downto -14);
Signal SumNode_Float416Output_1870: float (5 downto -14);
Signal ProductNode_Float1454Output_1871: float (5 downto -14);
Signal ProductNode_Float1455weight : float ( 5 downto -14 ) := to_float (0.870239,5,14);

Signal ProductNode_Float1455Output_1872: float (5 downto -14);
Signal SumNode_Float417Output_1873: float (5 downto -14);
Signal ProductNode_Float1456Output_1874: float (5 downto -14);
Signal ProductNode_Float1457weight : float ( 5 downto -14 ) := to_float (0.756327,5,14);

Signal ProductNode_Float1457Output_1875: float (5 downto -14);
Signal ProductNode_Float1458weight : float ( 5 downto -14 ) := to_float (0.890735,5,14);

Signal ProductNode_Float1458Output_1876: float (5 downto -14);
Signal ProductNode_Float1459weight : float ( 5 downto -14 ) := to_float (0.689002,5,14);

Signal ProductNode_Float1459Output_1877: float (5 downto -14);
Signal ProductNode_Float1460weight : float ( 5 downto -14 ) := to_float (0.966814,5,14);

Signal ProductNode_Float1460Output_1878: float (5 downto -14);
Signal SumNode_Float418Output_1879: float (5 downto -14);
Signal ProductNode_Float1461Output_1880: float (5 downto -14);
Signal ProductNode_Float1462weight : float ( 5 downto -14 ) := to_float (0.551341,5,14);

Signal ProductNode_Float1462Output_1881: float (5 downto -14);
Signal ProductNode_Float1463weight : float ( 5 downto -14 ) := to_float (0.795357,5,14);

Signal ProductNode_Float1463Output_1882: float (5 downto -14);
Signal ProductNode_Float1464weight : float ( 5 downto -14 ) := to_float (0.746308,5,14);

Signal ProductNode_Float1464Output_1883: float (5 downto -14);
Signal ProductNode_Float1465weight : float ( 5 downto -14 ) := to_float (0.989597,5,14);

Signal ProductNode_Float1465Output_1884: float (5 downto -14);
Signal ProductNode_Float1466weight : float ( 5 downto -14 ) := to_float (0.577708,5,14);

Signal ProductNode_Float1466Output_1885: float (5 downto -14);
Signal ProductNode_Float1467weight : float ( 5 downto -14 ) := to_float (0.618274,5,14);

Signal ProductNode_Float1467Output_1886: float (5 downto -14);
Signal SumNode_Float419Output_1887: float (5 downto -14);
Signal ProductNode_Float1468Output_1888: float (5 downto -14);
Signal ProductNode_Float1469weight : float ( 5 downto -14 ) := to_float (0.952809,5,14);

Signal ProductNode_Float1469Output_1889: float (5 downto -14);
Signal ProductNode_Float1470weight : float ( 5 downto -14 ) := to_float (0.495915,5,14);

Signal ProductNode_Float1470Output_1890: float (5 downto -14);
Signal ProductNode_Float1471weight : float ( 5 downto -14 ) := to_float (0.993928,5,14);

Signal ProductNode_Float1471Output_1891: float (5 downto -14);
Signal SumNode_Float420Output_1892: float (5 downto -14);
Signal ProductNode_Float1472Output_1893: float (5 downto -14);
Signal ProductNode_Float1473weight : float ( 5 downto -14 ) := to_float (0.551341,5,14);

Signal ProductNode_Float1473Output_1894: float (5 downto -14);
Signal ProductNode_Float1474weight : float ( 5 downto -14 ) := to_float (0.926235,5,14);

Signal ProductNode_Float1474Output_1895: float (5 downto -14);
Signal ProductNode_Float1475weight : float ( 5 downto -14 ) := to_float (0.616494,5,14);

Signal ProductNode_Float1475Output_1896: float (5 downto -14);
Signal ProductNode_Float1476weight : float ( 5 downto -14 ) := to_float (0.989597,5,14);

Signal ProductNode_Float1476Output_1897: float (5 downto -14);
Signal ProductNode_Float1477weight : float ( 5 downto -14 ) := to_float (0.986786,5,14);

Signal ProductNode_Float1477Output_1898: float (5 downto -14);
Signal ProductNode_Float1478weight : float ( 5 downto -14 ) := to_float (0.464416,5,14);

Signal ProductNode_Float1478Output_1899: float (5 downto -14);
Signal SumNode_Float421Output_1900: float (5 downto -14);
Signal ProductNode_Float1479Output_1901: float (5 downto -14);
Signal ProductNode_Float1480weight : float ( 5 downto -14 ) := to_float (0.770987,5,14);

Signal ProductNode_Float1480Output_1902: float (5 downto -14);
Signal SumNode_Float422Output_1903: float (5 downto -14);
Signal ProductNode_Float1481Output_1904: float (5 downto -14);
Signal ProductNode_Float1482weight : float ( 5 downto -14 ) := to_float (0.906302,5,14);

Signal ProductNode_Float1482Output_1905: float (5 downto -14);
Signal SumNode_Float423Output_1906: float (5 downto -14);
Signal ProductNode_Float1483Output_1907: float (5 downto -14);
Signal ProductNode_Float1484weight : float ( 5 downto -14 ) := to_float (0.923601,5,14);

Signal ProductNode_Float1484Output_1908: float (5 downto -14);
Signal ProductNode_Float1485weight : float ( 5 downto -14 ) := to_float (0.848299,5,14);

Signal ProductNode_Float1485Output_1909: float (5 downto -14);
Signal ProductNode_Float1486weight : float ( 5 downto -14 ) := to_float (0.562709,5,14);

Signal ProductNode_Float1486Output_1910: float (5 downto -14);
Signal ProductNode_Float1487weight : float ( 5 downto -14 ) := to_float (0.988453,5,14);

Signal ProductNode_Float1487Output_1911: float (5 downto -14);
Signal SumNode_Float424Output_1912: float (5 downto -14);
Signal ProductNode_Float1488Output_1913: float (5 downto -14);
Signal ProductNode_Float1489weight : float ( 5 downto -14 ) := to_float (0.870697,5,14);

Signal ProductNode_Float1489Output_1914: float (5 downto -14);
Signal ProductNode_Float1490weight : float ( 5 downto -14 ) := to_float (0.945793,5,14);

Signal ProductNode_Float1490Output_1915: float (5 downto -14);
Signal ProductNode_Float1491weight : float ( 5 downto -14 ) := to_float (0.729204,5,14);

Signal ProductNode_Float1491Output_1916: float (5 downto -14);
Signal ProductNode_Float1492weight : float ( 5 downto -14 ) := to_float (0.870404,5,14);

Signal ProductNode_Float1492Output_1917: float (5 downto -14);
Signal ProductNode_Float1493weight : float ( 5 downto -14 ) := to_float (0.780732,5,14);

Signal ProductNode_Float1493Output_1918: float (5 downto -14);
Signal ProductNode_Float1494weight : float ( 5 downto -14 ) := to_float (0.917308,5,14);

Signal ProductNode_Float1494Output_1919: float (5 downto -14);
Signal SumNode_Float425Output_1920: float (5 downto -14);
Signal ProductNode_Float1495Output_1921: float (5 downto -14);
Signal ProductNode_Float1496weight : float ( 5 downto -14 ) := to_float (0.979033,5,14);

Signal ProductNode_Float1496Output_1922: float (5 downto -14);
Signal ProductNode_Float1497weight : float ( 5 downto -14 ) := to_float (0.453222,5,14);

Signal ProductNode_Float1497Output_1923: float (5 downto -14);
Signal ProductNode_Float1498weight : float ( 5 downto -14 ) := to_float (0.996146,5,14);

Signal ProductNode_Float1498Output_1924: float (5 downto -14);
Signal SumNode_Float426Output_1925: float (5 downto -14);
Signal ProductNode_Float1499Output_1926: float (5 downto -14);
Signal ProductNode_Float1500weight : float ( 5 downto -14 ) := to_float (0.870697,5,14);

Signal ProductNode_Float1500Output_1927: float (5 downto -14);
Signal ProductNode_Float1501weight : float ( 5 downto -14 ) := to_float (0.753690,5,14);

Signal ProductNode_Float1501Output_1928: float (5 downto -14);
Signal ProductNode_Float1502weight : float ( 5 downto -14 ) := to_float (0.936763,5,14);

Signal ProductNode_Float1502Output_1929: float (5 downto -14);
Signal ProductNode_Float1503weight : float ( 5 downto -14 ) := to_float (0.870404,5,14);

Signal ProductNode_Float1503Output_1930: float (5 downto -14);
Signal ProductNode_Float1504weight : float ( 5 downto -14 ) := to_float (0.933776,5,14);

Signal ProductNode_Float1504Output_1931: float (5 downto -14);
Signal ProductNode_Float1505weight : float ( 5 downto -14 ) := to_float (0.973389,5,14);

Signal ProductNode_Float1505Output_1932: float (5 downto -14);
Signal SumNode_Float427Output_1933: float (5 downto -14);
Signal ProductNode_Float1506Output_1934: float (5 downto -14);
Signal ProductNode_Float1507weight : float ( 5 downto -14 ) := to_float (0.818419,5,14);

Signal ProductNode_Float1507Output_1935: float (5 downto -14);
Signal SumNode_Float428Output_1936: float (5 downto -14);
Signal ProductNode_Float1508Output_1937: float (5 downto -14);
Signal ProductNode_Float1509weight : float ( 5 downto -14 ) := to_float (0.940496,5,14);

Signal ProductNode_Float1509Output_1938: float (5 downto -14);
Signal ProductNode_Float1510weight : float ( 5 downto -14 ) := to_float (0.890735,5,14);

Signal ProductNode_Float1510Output_1939: float (5 downto -14);
Signal ProductNode_Float1511weight : float ( 5 downto -14 ) := to_float (0.382644,5,14);

Signal ProductNode_Float1511Output_1940: float (5 downto -14);
Signal ProductNode_Float1512weight : float ( 5 downto -14 ) := to_float (0.998354,5,14);

Signal ProductNode_Float1512Output_1941: float (5 downto -14);
Signal SumNode_Float429Output_1942: float (5 downto -14);
Signal ProductNode_Float1513Output_1943: float (5 downto -14);
Signal ProductNode_Float1514weight : float ( 5 downto -14 ) := to_float (0.551341,5,14);

Signal ProductNode_Float1514Output_1944: float (5 downto -14);
Signal ProductNode_Float1515weight : float ( 5 downto -14 ) := to_float (0.795357,5,14);

Signal ProductNode_Float1515Output_1945: float (5 downto -14);
Signal ProductNode_Float1516weight : float ( 5 downto -14 ) := to_float (0.948695,5,14);

Signal ProductNode_Float1516Output_1946: float (5 downto -14);
Signal ProductNode_Float1517weight : float ( 5 downto -14 ) := to_float (0.989597,5,14);

Signal ProductNode_Float1517Output_1947: float (5 downto -14);
Signal ProductNode_Float1518weight : float ( 5 downto -14 ) := to_float (0.577708,5,14);

Signal ProductNode_Float1518Output_1948: float (5 downto -14);
Signal ProductNode_Float1519weight : float ( 5 downto -14 ) := to_float (0.981240,5,14);

Signal ProductNode_Float1519Output_1949: float (5 downto -14);
Signal SumNode_Float430Output_1950: float (5 downto -14);
Signal ProductNode_Float1520Output_1951: float (5 downto -14);
Signal ProductNode_Float1521weight : float ( 5 downto -14 ) := to_float (0.960334,5,14);

Signal ProductNode_Float1521Output_1952: float (5 downto -14);
Signal ProductNode_Float1522weight : float ( 5 downto -14 ) := to_float (0.336149,5,14);

Signal ProductNode_Float1522Output_1953: float (5 downto -14);
Signal ProductNode_Float1523weight : float ( 5 downto -14 ) := to_float (0.999140,5,14);

Signal ProductNode_Float1523Output_1954: float (5 downto -14);
Signal SumNode_Float431Output_1955: float (5 downto -14);
Signal ProductNode_Float1524Output_1956: float (5 downto -14);
Signal ProductNode_Float1525weight : float ( 5 downto -14 ) := to_float (0.551341,5,14);

Signal ProductNode_Float1525Output_1957: float (5 downto -14);
Signal ProductNode_Float1526weight : float ( 5 downto -14 ) := to_float (0.926235,5,14);

Signal ProductNode_Float1526Output_1958: float (5 downto -14);
Signal ProductNode_Float1527weight : float ( 5 downto -14 ) := to_float (0.981519,5,14);

Signal ProductNode_Float1527Output_1959: float (5 downto -14);
Signal ProductNode_Float1528weight : float ( 5 downto -14 ) := to_float (0.989597,5,14);

Signal ProductNode_Float1528Output_1960: float (5 downto -14);
Signal ProductNode_Float1529weight : float ( 5 downto -14 ) := to_float (0.986786,5,14);

Signal ProductNode_Float1529Output_1961: float (5 downto -14);
Signal ProductNode_Float1530weight : float ( 5 downto -14 ) := to_float (0.995641,5,14);

Signal ProductNode_Float1530Output_1962: float (5 downto -14);
Signal SumNode_Float432Output_1963: float (5 downto -14);
Signal ProductNode_Float1531Output_1964: float (5 downto -14);
Signal ProductNode_Float1532weight : float ( 5 downto -14 ) := to_float (0.664315,5,14);

Signal ProductNode_Float1532Output_1965: float (5 downto -14);
Signal SumNode_Float433Output_1966: float (5 downto -14);
Signal ProductNode_Float1533Output_1967: float (5 downto -14);
Signal ProductNode_Float1534weight : float ( 5 downto -14 ) := to_float (0.978597,5,14);

Signal ProductNode_Float1534Output_1968: float (5 downto -14);
Signal SumNode_Float434Output_1969: float (5 downto -14);
Signal ProductNode_Float1535Output_1970: float (5 downto -14);
Signal ProductNode_Float1536weight : float ( 5 downto -14 ) := to_float (0.974456,5,14);

Signal ProductNode_Float1536Output_1971: float (5 downto -14);
Signal SumNode_Float435Output_1972: float (5 downto -14);
Signal ProductNode_Float1537Output_1973: float (5 downto -14);
Signal ProductNode_Float1538weight : float ( 5 downto -14 ) := to_float (0.970921,5,14);

Signal ProductNode_Float1538Output_1974: float (5 downto -14);
Signal ProductNode_Float1539weight : float ( 5 downto -14 ) := to_float (0.672140,5,14);

Signal ProductNode_Float1539Output_1975: float (5 downto -14);
Signal SumNode_Float436Output_1976: float (5 downto -14);
Signal ProductNode_Float1540Output_1977: float (5 downto -14);
Signal ProductNode_Float1541weight : float ( 5 downto -14 ) := to_float (0.989270,5,14);

Signal ProductNode_Float1541Output_1978: float (5 downto -14);
Signal ProductNode_Float1542weight : float ( 5 downto -14 ) := to_float (0.997554,5,14);

Signal ProductNode_Float1542Output_1979: float (5 downto -14);
Signal ProductNode_Float1543weight : float ( 5 downto -14 ) := to_float (0.414069,5,14);

Signal ProductNode_Float1543Output_1980: float (5 downto -14);
Signal SumNode_Float437Output_1981: float (5 downto -14);
Signal ProductNode_Float1544Output_1982: float (5 downto -14);
Signal ProductNode_Float1545weight : float ( 5 downto -14 ) := to_float (0.853307,5,14);

Signal ProductNode_Float1545Output_1983: float (5 downto -14);
Signal ProductNode_Float1546weight : float ( 5 downto -14 ) := to_float (0.886527,5,14);

Signal ProductNode_Float1546Output_1984: float (5 downto -14);
Signal SumNode_Float438Output_1985: float (5 downto -14);
Signal ProductNode_Float1547Output_1986: float (5 downto -14);
Signal ProductNode_Float1548weight : float ( 5 downto -14 ) := to_float (0.554692,5,14);

Signal ProductNode_Float1548Output_1987: float (5 downto -14);
Signal ProductNode_Float1549weight : float ( 5 downto -14 ) := to_float (0.989739,5,14);

Signal ProductNode_Float1549Output_1988: float (5 downto -14);
Signal ProductNode_Float1550weight : float ( 5 downto -14 ) := to_float (0.549861,5,14);

Signal ProductNode_Float1550Output_1989: float (5 downto -14);
Signal SumNode_Float439Output_1990: float (5 downto -14);
Signal ProductNode_Float1551Output_1991: float (5 downto -14);
Signal SumNode_Float440Output_1992: float (5 downto -14);
Signal ProductNode_Float1552Output_1993: float (5 downto -14);
Signal ProductNode_Float1553weight : float ( 5 downto -14 ) := to_float (0.994862,5,14);

Signal ProductNode_Float1553Output_1994: float (5 downto -14);
Signal ProductNode_Float1554weight : float ( 5 downto -14 ) := to_float (0.817897,5,14);

Signal ProductNode_Float1554Output_1995: float (5 downto -14);
Signal ProductNode_Float1555weight : float ( 5 downto -14 ) := to_float (0.912886,5,14);

Signal ProductNode_Float1555Output_1996: float (5 downto -14);
Signal SumNode_Float441Output_1997: float (5 downto -14);
Signal ProductNode_Float1556Output_1998: float (5 downto -14);
Signal ProductNode_Float1557weight : float ( 5 downto -14 ) := to_float (0.976301,5,14);

Signal ProductNode_Float1557Output_1999: float (5 downto -14);
Signal ProductNode_Float1558weight : float ( 5 downto -14 ) := to_float (0.988880,5,14);

Signal ProductNode_Float1558Output_2000: float (5 downto -14);
Signal ProductNode_Float1559weight : float ( 5 downto -14 ) := to_float (0.558577,5,14);

Signal ProductNode_Float1559Output_2001: float (5 downto -14);
Signal SumNode_Float442Output_2002: float (5 downto -14);
Signal ProductNode_Float1560Output_2003: float (5 downto -14);
Signal ProductNode_Float1561weight : float ( 5 downto -14 ) := to_float (0.731617,5,14);

Signal ProductNode_Float1561Output_2004: float (5 downto -14);
Signal ProductNode_Float1562weight : float ( 5 downto -14 ) := to_float (0.954043,5,14);

Signal ProductNode_Float1562Output_2005: float (5 downto -14);
Signal SumNode_Float443Output_2006: float (5 downto -14);
Signal ProductNode_Float1563Output_2007: float (5 downto -14);
Signal ProductNode_Float1564weight : float ( 5 downto -14 ) := to_float (0.646579,5,14);

Signal ProductNode_Float1564Output_2008: float (5 downto -14);
Signal ProductNode_Float1565weight : float ( 5 downto -14 ) := to_float (0.985013,5,14);

Signal ProductNode_Float1565Output_2009: float (5 downto -14);
Signal ProductNode_Float1566weight : float ( 5 downto -14 ) := to_float (0.592017,5,14);

Signal ProductNode_Float1566Output_2010: float (5 downto -14);
Signal SumNode_Float444Output_2011: float (5 downto -14);
Signal ProductNode_Float1567Output_2012: float (5 downto -14);
Signal SumNode_Float445Output_2013: float (5 downto -14);
Signal ProductNode_Float1568Output_2014: float (5 downto -14);
Signal ProductNode_Float1569weight : float ( 5 downto -14 ) := to_float (0.479802,5,14);

Signal ProductNode_Float1569Output_2015: float (5 downto -14);
Signal SumNode_Float446Output_2016: float (5 downto -14);
Signal ProductNode_Float1570Output_2017: float (5 downto -14);
Signal ProductNode_Float1571weight : float ( 5 downto -14 ) := to_float (0.807423,5,14);

Signal ProductNode_Float1571Output_2018: float (5 downto -14);
Signal ProductNode_Float1572weight : float ( 5 downto -14 ) := to_float (0.919372,5,14);

Signal ProductNode_Float1572Output_2019: float (5 downto -14);
Signal SumNode_Float447Output_2020: float (5 downto -14);
Signal ProductNode_Float1573Output_2021: float (5 downto -14);
Signal ProductNode_Float1574weight : float ( 5 downto -14 ) := to_float (0.694473,5,14);

Signal ProductNode_Float1574Output_2022: float (5 downto -14);
Signal ProductNode_Float1575weight : float ( 5 downto -14 ) := to_float (0.843444,5,14);

Signal ProductNode_Float1575Output_2023: float (5 downto -14);
Signal ProductNode_Float1576weight : float ( 5 downto -14 ) := to_float (0.682797,5,14);

Signal ProductNode_Float1576Output_2024: float (5 downto -14);
Signal ProductNode_Float1577weight : float ( 5 downto -14 ) := to_float (0.968381,5,14);

Signal ProductNode_Float1577Output_2025: float (5 downto -14);
Signal SumNode_Float448Output_2026: float (5 downto -14);
Signal ProductNode_Float1578Output_2027: float (5 downto -14);
Signal ProductNode_Float1579weight : float ( 5 downto -14 ) := to_float (0.965376,5,14);

Signal ProductNode_Float1579Output_2028: float (5 downto -14);
Signal ProductNode_Float1580weight : float ( 5 downto -14 ) := to_float (0.697447,5,14);

Signal ProductNode_Float1580Output_2029: float (5 downto -14);
Signal SumNode_Float449Output_2030: float (5 downto -14);
Signal ProductNode_Float1581Output_2031: float (5 downto -14);
Signal ProductNode_Float1582weight : float ( 5 downto -14 ) := to_float (0.970921,5,14);

Signal ProductNode_Float1582Output_2032: float (5 downto -14);
Signal ProductNode_Float1583weight : float ( 5 downto -14 ) := to_float (0.672140,5,14);

Signal ProductNode_Float1583Output_2033: float (5 downto -14);
Signal SumNode_Float450Output_2034: float (5 downto -14);
Signal ProductNode_Float1584Output_2035: float (5 downto -14);
Signal ProductNode_Float1585weight : float ( 5 downto -14 ) := to_float (0.989270,5,14);

Signal ProductNode_Float1585Output_2036: float (5 downto -14);
Signal ProductNode_Float1586weight : float ( 5 downto -14 ) := to_float (0.997554,5,14);

Signal ProductNode_Float1586Output_2037: float (5 downto -14);
Signal ProductNode_Float1587weight : float ( 5 downto -14 ) := to_float (0.414069,5,14);

Signal ProductNode_Float1587Output_2038: float (5 downto -14);
Signal SumNode_Float451Output_2039: float (5 downto -14);
Signal ProductNode_Float1588Output_2040: float (5 downto -14);
Signal ProductNode_Float1589weight : float ( 5 downto -14 ) := to_float (0.853307,5,14);

Signal ProductNode_Float1589Output_2041: float (5 downto -14);
Signal ProductNode_Float1590weight : float ( 5 downto -14 ) := to_float (0.886527,5,14);

Signal ProductNode_Float1590Output_2042: float (5 downto -14);
Signal SumNode_Float452Output_2043: float (5 downto -14);
Signal ProductNode_Float1591Output_2044: float (5 downto -14);
Signal ProductNode_Float1592weight : float ( 5 downto -14 ) := to_float (0.554692,5,14);

Signal ProductNode_Float1592Output_2045: float (5 downto -14);
Signal ProductNode_Float1593weight : float ( 5 downto -14 ) := to_float (0.989739,5,14);

Signal ProductNode_Float1593Output_2046: float (5 downto -14);
Signal ProductNode_Float1594weight : float ( 5 downto -14 ) := to_float (0.549861,5,14);

Signal ProductNode_Float1594Output_2047: float (5 downto -14);
Signal SumNode_Float453Output_2048: float (5 downto -14);
Signal ProductNode_Float1595Output_2049: float (5 downto -14);
Signal SumNode_Float454Output_2050: float (5 downto -14);
Signal ProductNode_Float1596Output_2051: float (5 downto -14);
Signal ProductNode_Float1597weight : float ( 5 downto -14 ) := to_float (0.970629,5,14);

Signal ProductNode_Float1597Output_2052: float (5 downto -14);
Signal ProductNode_Float1598weight : float ( 5 downto -14 ) := to_float (0.817897,5,14);

Signal ProductNode_Float1598Output_2053: float (5 downto -14);
Signal ProductNode_Float1599weight : float ( 5 downto -14 ) := to_float (0.912886,5,14);

Signal ProductNode_Float1599Output_2054: float (5 downto -14);
Signal SumNode_Float455Output_2055: float (5 downto -14);
Signal ProductNode_Float1600Output_2056: float (5 downto -14);
Signal ProductNode_Float1601weight : float ( 5 downto -14 ) := to_float (0.976301,5,14);

Signal ProductNode_Float1601Output_2057: float (5 downto -14);
Signal ProductNode_Float1602weight : float ( 5 downto -14 ) := to_float (0.988880,5,14);

Signal ProductNode_Float1602Output_2058: float (5 downto -14);
Signal ProductNode_Float1603weight : float ( 5 downto -14 ) := to_float (0.558577,5,14);

Signal ProductNode_Float1603Output_2059: float (5 downto -14);
Signal SumNode_Float456Output_2060: float (5 downto -14);
Signal ProductNode_Float1604Output_2061: float (5 downto -14);
Signal ProductNode_Float1605weight : float ( 5 downto -14 ) := to_float (0.731617,5,14);

Signal ProductNode_Float1605Output_2062: float (5 downto -14);
Signal ProductNode_Float1606weight : float ( 5 downto -14 ) := to_float (0.954043,5,14);

Signal ProductNode_Float1606Output_2063: float (5 downto -14);
Signal SumNode_Float457Output_2064: float (5 downto -14);
Signal ProductNode_Float1607Output_2065: float (5 downto -14);
Signal ProductNode_Float1608weight : float ( 5 downto -14 ) := to_float (0.646579,5,14);

Signal ProductNode_Float1608Output_2066: float (5 downto -14);
Signal ProductNode_Float1609weight : float ( 5 downto -14 ) := to_float (0.985013,5,14);

Signal ProductNode_Float1609Output_2067: float (5 downto -14);
Signal ProductNode_Float1610weight : float ( 5 downto -14 ) := to_float (0.592017,5,14);

Signal ProductNode_Float1610Output_2068: float (5 downto -14);
Signal SumNode_Float458Output_2069: float (5 downto -14);
Signal ProductNode_Float1611Output_2070: float (5 downto -14);
Signal SumNode_Float459Output_2071: float (5 downto -14);
Signal ProductNode_Float1612Output_2072: float (5 downto -14);
Signal ProductNode_Float1613weight : float ( 5 downto -14 ) := to_float (0.673404,5,14);

Signal ProductNode_Float1613Output_2073: float (5 downto -14);
Signal SumNode_Float460Output_2074: float (5 downto -14);
Signal ProductNode_Float1614Output_2075: float (5 downto -14);
Signal ProductNode_Float1615weight : float ( 5 downto -14 ) := to_float (0.623360,5,14);

Signal ProductNode_Float1615Output_2076: float (5 downto -14);
Signal ProductNode_Float1616weight : float ( 5 downto -14 ) := to_float (0.980424,5,14);

Signal ProductNode_Float1616Output_2077: float (5 downto -14);
Signal SumNode_Float461Output_2078: float (5 downto -14);
Signal ProductNode_Float1617Output_2079: float (5 downto -14);
Signal ProductNode_Float1618weight : float ( 5 downto -14 ) := to_float (0.694473,5,14);

Signal ProductNode_Float1618Output_2080: float (5 downto -14);
Signal ProductNode_Float1619weight : float ( 5 downto -14 ) := to_float (0.894649,5,14);

Signal ProductNode_Float1619Output_2081: float (5 downto -14);
Signal ProductNode_Float1620weight : float ( 5 downto -14 ) := to_float (0.482891,5,14);

Signal ProductNode_Float1620Output_2082: float (5 downto -14);
Signal ProductNode_Float1621weight : float ( 5 downto -14 ) := to_float (0.994693,5,14);

Signal ProductNode_Float1621Output_2083: float (5 downto -14);
Signal SumNode_Float462Output_2084: float (5 downto -14);
Signal ProductNode_Float1622Output_2085: float (5 downto -14);
Signal ProductNode_Float1623weight : float ( 5 downto -14 ) := to_float (0.965376,5,14);

Signal ProductNode_Float1623Output_2086: float (5 downto -14);
Signal ProductNode_Float1624weight : float ( 5 downto -14 ) := to_float (0.964572,5,14);

Signal ProductNode_Float1624Output_2087: float (5 downto -14);
Signal SumNode_Float463Output_2088: float (5 downto -14);
Signal ProductNode_Float1625Output_2089: float (5 downto -14);
Signal SumNode_Float464Output_2090: float (5 downto -14);
Signal ProductNode_Float1626Output_2091: float (5 downto -14);
Signal ProductNode_Float1627weight : float ( 5 downto -14 ) := to_float (0.768486,5,14);

Signal ProductNode_Float1627Output_2092: float (5 downto -14);
Signal ProductNode_Float1628weight : float ( 5 downto -14 ) := to_float (0.970921,5,14);

Signal ProductNode_Float1628Output_2093: float (5 downto -14);
Signal ProductNode_Float1629weight : float ( 5 downto -14 ) := to_float (0.672140,5,14);

Signal ProductNode_Float1629Output_2094: float (5 downto -14);
Signal SumNode_Float465Output_2095: float (5 downto -14);
Signal ProductNode_Float1630Output_2096: float (5 downto -14);
Signal ProductNode_Float1631weight : float ( 5 downto -14 ) := to_float (0.989270,5,14);

Signal ProductNode_Float1631Output_2097: float (5 downto -14);
Signal ProductNode_Float1632weight : float ( 5 downto -14 ) := to_float (0.966381,5,14);

Signal ProductNode_Float1632Output_2098: float (5 downto -14);
Signal ProductNode_Float1633weight : float ( 5 downto -14 ) := to_float (0.690672,5,14);

Signal ProductNode_Float1633Output_2099: float (5 downto -14);
Signal SumNode_Float466Output_2100: float (5 downto -14);
Signal ProductNode_Float1634Output_2101: float (5 downto -14);
Signal ProductNode_Float1635weight : float ( 5 downto -14 ) := to_float (0.853307,5,14);

Signal ProductNode_Float1635Output_2102: float (5 downto -14);
Signal ProductNode_Float1636weight : float ( 5 downto -14 ) := to_float (0.886527,5,14);

Signal ProductNode_Float1636Output_2103: float (5 downto -14);
Signal SumNode_Float467Output_2104: float (5 downto -14);
Signal ProductNode_Float1637Output_2105: float (5 downto -14);
Signal ProductNode_Float1638weight : float ( 5 downto -14 ) := to_float (0.554692,5,14);

Signal ProductNode_Float1638Output_2106: float (5 downto -14);
Signal ProductNode_Float1639weight : float ( 5 downto -14 ) := to_float (0.941870,5,14);

Signal ProductNode_Float1639Output_2107: float (5 downto -14);
Signal ProductNode_Float1640weight : float ( 5 downto -14 ) := to_float (0.763101,5,14);

Signal ProductNode_Float1640Output_2108: float (5 downto -14);
Signal SumNode_Float468Output_2109: float (5 downto -14);
Signal ProductNode_Float1641Output_2110: float (5 downto -14);
Signal SumNode_Float469Output_2111: float (5 downto -14);
Signal ProductNode_Float1642Output_2112: float (5 downto -14);
Signal ProductNode_Float1643weight : float ( 5 downto -14 ) := to_float (0.951966,5,14);

Signal ProductNode_Float1643Output_2113: float (5 downto -14);
Signal ProductNode_Float1644weight : float ( 5 downto -14 ) := to_float (0.817897,5,14);

Signal ProductNode_Float1644Output_2114: float (5 downto -14);
Signal ProductNode_Float1645weight : float ( 5 downto -14 ) := to_float (0.912886,5,14);

Signal ProductNode_Float1645Output_2115: float (5 downto -14);
Signal SumNode_Float470Output_2116: float (5 downto -14);
Signal ProductNode_Float1646Output_2117: float (5 downto -14);
Signal ProductNode_Float1647weight : float ( 5 downto -14 ) := to_float (0.976301,5,14);

Signal ProductNode_Float1647Output_2118: float (5 downto -14);
Signal ProductNode_Float1648weight : float ( 5 downto -14 ) := to_float (0.909585,5,14);

Signal ProductNode_Float1648Output_2119: float (5 downto -14);
Signal ProductNode_Float1649weight : float ( 5 downto -14 ) := to_float (0.822920,5,14);

Signal ProductNode_Float1649Output_2120: float (5 downto -14);
Signal SumNode_Float471Output_2121: float (5 downto -14);
Signal ProductNode_Float1650Output_2122: float (5 downto -14);
Signal ProductNode_Float1651weight : float ( 5 downto -14 ) := to_float (0.731617,5,14);

Signal ProductNode_Float1651Output_2123: float (5 downto -14);
Signal ProductNode_Float1652weight : float ( 5 downto -14 ) := to_float (0.954043,5,14);

Signal ProductNode_Float1652Output_2124: float (5 downto -14);
Signal SumNode_Float472Output_2125: float (5 downto -14);
Signal ProductNode_Float1653Output_2126: float (5 downto -14);
Signal ProductNode_Float1654weight : float ( 5 downto -14 ) := to_float (0.646579,5,14);

Signal ProductNode_Float1654Output_2127: float (5 downto -14);
Signal ProductNode_Float1655weight : float ( 5 downto -14 ) := to_float (0.790147,5,14);

Signal ProductNode_Float1655Output_2128: float (5 downto -14);
Signal ProductNode_Float1656weight : float ( 5 downto -14 ) := to_float (0.929014,5,14);

Signal ProductNode_Float1656Output_2129: float (5 downto -14);
Signal SumNode_Float473Output_2130: float (5 downto -14);
Signal ProductNode_Float1657Output_2131: float (5 downto -14);
Signal SumNode_Float474Output_2132: float (5 downto -14);
Signal ProductNode_Float1658Output_2133: float (5 downto -14);
Signal ProductNode_Float1659weight : float ( 5 downto -14 ) := to_float (0.737500,5,14);

Signal ProductNode_Float1659Output_2134: float (5 downto -14);
Signal SumNode_Float475Output_2135: float (5 downto -14);
Signal ProductNode_Float1660Output_2136: float (5 downto -14);
Signal ProductNode_Float1661weight : float ( 5 downto -14 ) := to_float (0.807423,5,14);

Signal ProductNode_Float1661Output_2137: float (5 downto -14);
Signal ProductNode_Float1662weight : float ( 5 downto -14 ) := to_float (0.919372,5,14);

Signal ProductNode_Float1662Output_2138: float (5 downto -14);
Signal SumNode_Float476Output_2139: float (5 downto -14);
Signal ProductNode_Float1663Output_2140: float (5 downto -14);
Signal ProductNode_Float1664weight : float ( 5 downto -14 ) := to_float (0.579487,5,14);

Signal ProductNode_Float1664Output_2141: float (5 downto -14);
Signal ProductNode_Float1665weight : float ( 5 downto -14 ) := to_float (0.790558,5,14);

Signal ProductNode_Float1665Output_2142: float (5 downto -14);
Signal ProductNode_Float1666weight : float ( 5 downto -14 ) := to_float (0.682797,5,14);

Signal ProductNode_Float1666Output_2143: float (5 downto -14);
Signal ProductNode_Float1667weight : float ( 5 downto -14 ) := to_float (0.968381,5,14);

Signal ProductNode_Float1667Output_2144: float (5 downto -14);
Signal SumNode_Float477Output_2145: float (5 downto -14);
Signal ProductNode_Float1668Output_2146: float (5 downto -14);
Signal ProductNode_Float1669weight : float ( 5 downto -14 ) := to_float (0.986575,5,14);

Signal ProductNode_Float1669Output_2147: float (5 downto -14);
Signal ProductNode_Float1670weight : float ( 5 downto -14 ) := to_float (0.578242,5,14);

Signal ProductNode_Float1670Output_2148: float (5 downto -14);
Signal SumNode_Float478Output_2149: float (5 downto -14);
Signal ProductNode_Float1671Output_2150: float (5 downto -14);
Signal ProductNode_Float1672weight : float ( 5 downto -14 ) := to_float (0.970921,5,14);

Signal ProductNode_Float1672Output_2151: float (5 downto -14);
Signal ProductNode_Float1673weight : float ( 5 downto -14 ) := to_float (0.672140,5,14);

Signal ProductNode_Float1673Output_2152: float (5 downto -14);
Signal SumNode_Float479Output_2153: float (5 downto -14);
Signal ProductNode_Float1674Output_2154: float (5 downto -14);
Signal ProductNode_Float1675weight : float ( 5 downto -14 ) := to_float (0.989270,5,14);

Signal ProductNode_Float1675Output_2155: float (5 downto -14);
Signal ProductNode_Float1676weight : float ( 5 downto -14 ) := to_float (0.966381,5,14);

Signal ProductNode_Float1676Output_2156: float (5 downto -14);
Signal ProductNode_Float1677weight : float ( 5 downto -14 ) := to_float (0.690672,5,14);

Signal ProductNode_Float1677Output_2157: float (5 downto -14);
Signal SumNode_Float480Output_2158: float (5 downto -14);
Signal ProductNode_Float1678Output_2159: float (5 downto -14);
Signal ProductNode_Float1679weight : float ( 5 downto -14 ) := to_float (0.853307,5,14);

Signal ProductNode_Float1679Output_2160: float (5 downto -14);
Signal ProductNode_Float1680weight : float ( 5 downto -14 ) := to_float (0.886527,5,14);

Signal ProductNode_Float1680Output_2161: float (5 downto -14);
Signal SumNode_Float481Output_2162: float (5 downto -14);
Signal ProductNode_Float1681Output_2163: float (5 downto -14);
Signal ProductNode_Float1682weight : float ( 5 downto -14 ) := to_float (0.554692,5,14);

Signal ProductNode_Float1682Output_2164: float (5 downto -14);
Signal ProductNode_Float1683weight : float ( 5 downto -14 ) := to_float (0.941870,5,14);

Signal ProductNode_Float1683Output_2165: float (5 downto -14);
Signal ProductNode_Float1684weight : float ( 5 downto -14 ) := to_float (0.763101,5,14);

Signal ProductNode_Float1684Output_2166: float (5 downto -14);
Signal SumNode_Float482Output_2167: float (5 downto -14);
Signal ProductNode_Float1685Output_2168: float (5 downto -14);
Signal SumNode_Float483Output_2169: float (5 downto -14);
Signal ProductNode_Float1686Output_2170: float (5 downto -14);
Signal ProductNode_Float1687weight : float ( 5 downto -14 ) := to_float (0.840616,5,14);

Signal ProductNode_Float1687Output_2171: float (5 downto -14);
Signal ProductNode_Float1688weight : float ( 5 downto -14 ) := to_float (0.817897,5,14);

Signal ProductNode_Float1688Output_2172: float (5 downto -14);
Signal ProductNode_Float1689weight : float ( 5 downto -14 ) := to_float (0.912886,5,14);

Signal ProductNode_Float1689Output_2173: float (5 downto -14);
Signal SumNode_Float484Output_2174: float (5 downto -14);
Signal ProductNode_Float1690Output_2175: float (5 downto -14);
Signal ProductNode_Float1691weight : float ( 5 downto -14 ) := to_float (0.976301,5,14);

Signal ProductNode_Float1691Output_2176: float (5 downto -14);
Signal ProductNode_Float1692weight : float ( 5 downto -14 ) := to_float (0.909585,5,14);

Signal ProductNode_Float1692Output_2177: float (5 downto -14);
Signal ProductNode_Float1693weight : float ( 5 downto -14 ) := to_float (0.822920,5,14);

Signal ProductNode_Float1693Output_2178: float (5 downto -14);
Signal SumNode_Float485Output_2179: float (5 downto -14);
Signal ProductNode_Float1694Output_2180: float (5 downto -14);
Signal ProductNode_Float1695weight : float ( 5 downto -14 ) := to_float (0.731617,5,14);

Signal ProductNode_Float1695Output_2181: float (5 downto -14);
Signal ProductNode_Float1696weight : float ( 5 downto -14 ) := to_float (0.954043,5,14);

Signal ProductNode_Float1696Output_2182: float (5 downto -14);
Signal SumNode_Float486Output_2183: float (5 downto -14);
Signal ProductNode_Float1697Output_2184: float (5 downto -14);
Signal ProductNode_Float1698weight : float ( 5 downto -14 ) := to_float (0.646579,5,14);

Signal ProductNode_Float1698Output_2185: float (5 downto -14);
Signal ProductNode_Float1699weight : float ( 5 downto -14 ) := to_float (0.790147,5,14);

Signal ProductNode_Float1699Output_2186: float (5 downto -14);
Signal ProductNode_Float1700weight : float ( 5 downto -14 ) := to_float (0.929014,5,14);

Signal ProductNode_Float1700Output_2187: float (5 downto -14);
Signal SumNode_Float487Output_2188: float (5 downto -14);
Signal ProductNode_Float1701Output_2189: float (5 downto -14);
Signal SumNode_Float488Output_2190: float (5 downto -14);
Signal ProductNode_Float1702Output_2191: float (5 downto -14);
Signal ProductNode_Float1703weight : float ( 5 downto -14 ) := to_float (0.896858,5,14);

Signal ProductNode_Float1703Output_2192: float (5 downto -14);
Signal SumNode_Float489Output_2193: float (5 downto -14);
Signal ProductNode_Float1704Output_2194: float (5 downto -14);
Signal ProductNode_Float1705weight : float ( 5 downto -14 ) := to_float (0.623360,5,14);

Signal ProductNode_Float1705Output_2195: float (5 downto -14);
Signal ProductNode_Float1706weight : float ( 5 downto -14 ) := to_float (0.980424,5,14);

Signal ProductNode_Float1706Output_2196: float (5 downto -14);
Signal SumNode_Float490Output_2197: float (5 downto -14);
Signal ProductNode_Float1707Output_2198: float (5 downto -14);
Signal ProductNode_Float1708weight : float ( 5 downto -14 ) := to_float (0.579487,5,14);

Signal ProductNode_Float1708Output_2199: float (5 downto -14);
Signal ProductNode_Float1709weight : float ( 5 downto -14 ) := to_float (0.928799,5,14);

Signal ProductNode_Float1709Output_2200: float (5 downto -14);
Signal ProductNode_Float1710weight : float ( 5 downto -14 ) := to_float (0.482891,5,14);

Signal ProductNode_Float1710Output_2201: float (5 downto -14);
Signal ProductNode_Float1711weight : float ( 5 downto -14 ) := to_float (0.994693,5,14);

Signal ProductNode_Float1711Output_2202: float (5 downto -14);
Signal SumNode_Float491Output_2203: float (5 downto -14);
Signal ProductNode_Float1712Output_2204: float (5 downto -14);
Signal ProductNode_Float1713weight : float ( 5 downto -14 ) := to_float (0.986575,5,14);

Signal ProductNode_Float1713Output_2205: float (5 downto -14);
Signal ProductNode_Float1714weight : float ( 5 downto -14 ) := to_float (0.986723,5,14);

Signal ProductNode_Float1714Output_2206: float (5 downto -14);
Signal SumNode_Float492Output_2207: float (5 downto -14);
Signal ProductNode_Float1715Output_2208: float (5 downto -14);
Signal SumNode_Float493Output_2209: float (5 downto -14);
Signal ProductNode_Float1716Output_2210: float (5 downto -14);
Signal ProductNode_Float1717weight : float ( 5 downto -14 ) := to_float (0.939505,5,14);

Signal ProductNode_Float1717Output_2211: float (5 downto -14);
Signal SumNode_Float494Output_2212: float (5 downto -14);
Signal ProductNode_Float1718Output_2213: float (5 downto -14);
Signal SumNode_Float495Output_2214: float (5 downto -14);
Signal ProductNode_Float1719Output_2215: float (5 downto -14);
Signal ProductNode_Float1720weight : float ( 5 downto -14 ) := to_float (0.848299,5,14);

Signal ProductNode_Float1720Output_2216: float (5 downto -14);
Signal ProductNode_Float1721weight : float ( 5 downto -14 ) := to_float (0.895308,5,14);

Signal ProductNode_Float1721Output_2217: float (5 downto -14);
Signal ProductNode_Float1722weight : float ( 5 downto -14 ) := to_float (0.842608,5,14);

Signal ProductNode_Float1722Output_2218: float (5 downto -14);
Signal SumNode_Float496Output_2219: float (5 downto -14);
Signal ProductNode_Float1723Output_2220: float (5 downto -14);
Signal ProductNode_Float1724weight : float ( 5 downto -14 ) := to_float (0.870697,5,14);

Signal ProductNode_Float1724Output_2221: float (5 downto -14);
Signal ProductNode_Float1725weight : float ( 5 downto -14 ) := to_float (0.945793,5,14);

Signal ProductNode_Float1725Output_2222: float (5 downto -14);
Signal ProductNode_Float1726weight : float ( 5 downto -14 ) := to_float (0.954870,5,14);

Signal ProductNode_Float1726Output_2223: float (5 downto -14);
Signal ProductNode_Float1727weight : float ( 5 downto -14 ) := to_float (0.870404,5,14);

Signal ProductNode_Float1727Output_2224: float (5 downto -14);
Signal ProductNode_Float1728weight : float ( 5 downto -14 ) := to_float (0.780732,5,14);

Signal ProductNode_Float1728Output_2225: float (5 downto -14);
Signal ProductNode_Float1729weight : float ( 5 downto -14 ) := to_float (0.810846,5,14);

Signal ProductNode_Float1729Output_2226: float (5 downto -14);
Signal SumNode_Float497Output_2227: float (5 downto -14);
Signal ProductNode_Float1730Output_2228: float (5 downto -14);
Signal ProductNode_Float1731weight : float ( 5 downto -14 ) := to_float (0.531606,5,14);

Signal ProductNode_Float1731Output_2229: float (5 downto -14);
Signal ProductNode_Float1732weight : float ( 5 downto -14 ) := to_float (0.669241,5,14);

Signal ProductNode_Float1732Output_2230: float (5 downto -14);
Signal ProductNode_Float1733weight : float ( 5 downto -14 ) := to_float (0.971580,5,14);

Signal ProductNode_Float1733Output_2231: float (5 downto -14);
Signal SumNode_Float498Output_2232: float (5 downto -14);
Signal ProductNode_Float1734Output_2233: float (5 downto -14);
Signal ProductNode_Float1735weight : float ( 5 downto -14 ) := to_float (0.870697,5,14);

Signal ProductNode_Float1735Output_2234: float (5 downto -14);
Signal ProductNode_Float1736weight : float ( 5 downto -14 ) := to_float (0.753690,5,14);

Signal ProductNode_Float1736Output_2235: float (5 downto -14);
Signal ProductNode_Float1737weight : float ( 5 downto -14 ) := to_float (0.774480,5,14);

Signal ProductNode_Float1737Output_2236: float (5 downto -14);
Signal ProductNode_Float1738weight : float ( 5 downto -14 ) := to_float (0.870404,5,14);

Signal ProductNode_Float1738Output_2237: float (5 downto -14);
Signal ProductNode_Float1739weight : float ( 5 downto -14 ) := to_float (0.933776,5,14);

Signal ProductNode_Float1739Output_2238: float (5 downto -14);
Signal ProductNode_Float1740weight : float ( 5 downto -14 ) := to_float (0.660973,5,14);

Signal ProductNode_Float1740Output_2239: float (5 downto -14);
Signal SumNode_Float499Output_2240: float (5 downto -14);
Signal ProductNode_Float1741Output_2241: float (5 downto -14);
Signal ProductNode_Float1742weight : float ( 5 downto -14 ) := to_float (0.870862,5,14);

Signal ProductNode_Float1742Output_2242: float (5 downto -14);
Signal SumNode_Float500Output_2243: float (5 downto -14);
Signal ProductNode_Float1743Output_2244: float (5 downto -14);
Signal ProductNode_Float1744weight : float ( 5 downto -14 ) := to_float (0.850730,5,14);

Signal ProductNode_Float1744Output_2245: float (5 downto -14);
Signal ProductNode_Float1745weight : float ( 5 downto -14 ) := to_float (0.890735,5,14);

Signal ProductNode_Float1745Output_2246: float (5 downto -14);
Signal ProductNode_Float1746weight : float ( 5 downto -14 ) := to_float (0.689002,5,14);

Signal ProductNode_Float1746Output_2247: float (5 downto -14);
Signal ProductNode_Float1747weight : float ( 5 downto -14 ) := to_float (0.966814,5,14);

Signal ProductNode_Float1747Output_2248: float (5 downto -14);
Signal SumNode_Float501Output_2249: float (5 downto -14);
Signal ProductNode_Float1748Output_2250: float (5 downto -14);
Signal ProductNode_Float1749weight : float ( 5 downto -14 ) := to_float (0.551341,5,14);

Signal ProductNode_Float1749Output_2251: float (5 downto -14);
Signal ProductNode_Float1750weight : float ( 5 downto -14 ) := to_float (0.795357,5,14);

Signal ProductNode_Float1750Output_2252: float (5 downto -14);
Signal ProductNode_Float1751weight : float ( 5 downto -14 ) := to_float (0.746308,5,14);

Signal ProductNode_Float1751Output_2253: float (5 downto -14);
Signal ProductNode_Float1752weight : float ( 5 downto -14 ) := to_float (0.989597,5,14);

Signal ProductNode_Float1752Output_2254: float (5 downto -14);
Signal ProductNode_Float1753weight : float ( 5 downto -14 ) := to_float (0.577708,5,14);

Signal ProductNode_Float1753Output_2255: float (5 downto -14);
Signal ProductNode_Float1754weight : float ( 5 downto -14 ) := to_float (0.618274,5,14);

Signal ProductNode_Float1754Output_2256: float (5 downto -14);
Signal SumNode_Float502Output_2257: float (5 downto -14);
Signal ProductNode_Float1755Output_2258: float (5 downto -14);
Signal ProductNode_Float1756weight : float ( 5 downto -14 ) := to_float (0.735141,5,14);

Signal ProductNode_Float1756Output_2259: float (5 downto -14);
Signal ProductNode_Float1757weight : float ( 5 downto -14 ) := to_float (0.495915,5,14);

Signal ProductNode_Float1757Output_2260: float (5 downto -14);
Signal ProductNode_Float1758weight : float ( 5 downto -14 ) := to_float (0.993928,5,14);

Signal ProductNode_Float1758Output_2261: float (5 downto -14);
Signal SumNode_Float503Output_2262: float (5 downto -14);
Signal ProductNode_Float1759Output_2263: float (5 downto -14);
Signal ProductNode_Float1760weight : float ( 5 downto -14 ) := to_float (0.551341,5,14);

Signal ProductNode_Float1760Output_2264: float (5 downto -14);
Signal ProductNode_Float1761weight : float ( 5 downto -14 ) := to_float (0.926235,5,14);

Signal ProductNode_Float1761Output_2265: float (5 downto -14);
Signal ProductNode_Float1762weight : float ( 5 downto -14 ) := to_float (0.616494,5,14);

Signal ProductNode_Float1762Output_2266: float (5 downto -14);
Signal ProductNode_Float1763weight : float ( 5 downto -14 ) := to_float (0.989597,5,14);

Signal ProductNode_Float1763Output_2267: float (5 downto -14);
Signal ProductNode_Float1764weight : float ( 5 downto -14 ) := to_float (0.986786,5,14);

Signal ProductNode_Float1764Output_2268: float (5 downto -14);
Signal ProductNode_Float1765weight : float ( 5 downto -14 ) := to_float (0.464416,5,14);

Signal ProductNode_Float1765Output_2269: float (5 downto -14);
Signal SumNode_Float504Output_2270: float (5 downto -14);
Signal ProductNode_Float1766Output_2271: float (5 downto -14);
Signal ProductNode_Float1767weight : float ( 5 downto -14 ) := to_float (0.938375,5,14);

Signal ProductNode_Float1767Output_2272: float (5 downto -14);
Signal SumNode_Float505Output_2273: float (5 downto -14);
Signal ProductNode_Float1768Output_2274: float (5 downto -14);
Signal ProductNode_Float1769weight : float ( 5 downto -14 ) := to_float (0.635106,5,14);

Signal ProductNode_Float1769Output_2275: float (5 downto -14);
Signal SumNode_Float506Output_2276: float (5 downto -14);
Signal ProductNode_Float1770Output_2277: float (5 downto -14);
Signal ProductNode_Float1771weight : float ( 5 downto -14 ) := to_float (0.677835,5,14);

Signal ProductNode_Float1771Output_2278: float (5 downto -14);
Signal ProductNode_Float1772weight : float ( 5 downto -14 ) := to_float (0.848299,5,14);

Signal ProductNode_Float1772Output_2279: float (5 downto -14);
Signal ProductNode_Float1773weight : float ( 5 downto -14 ) := to_float (0.562709,5,14);

Signal ProductNode_Float1773Output_2280: float (5 downto -14);
Signal ProductNode_Float1774weight : float ( 5 downto -14 ) := to_float (0.988453,5,14);

Signal ProductNode_Float1774Output_2281: float (5 downto -14);
Signal SumNode_Float507Output_2282: float (5 downto -14);
Signal ProductNode_Float1775Output_2283: float (5 downto -14);
Signal ProductNode_Float1776weight : float ( 5 downto -14 ) := to_float (0.870697,5,14);

Signal ProductNode_Float1776Output_2284: float (5 downto -14);
Signal ProductNode_Float1777weight : float ( 5 downto -14 ) := to_float (0.945793,5,14);

Signal ProductNode_Float1777Output_2285: float (5 downto -14);
Signal ProductNode_Float1778weight : float ( 5 downto -14 ) := to_float (0.729204,5,14);

Signal ProductNode_Float1778Output_2286: float (5 downto -14);
Signal ProductNode_Float1779weight : float ( 5 downto -14 ) := to_float (0.870404,5,14);

Signal ProductNode_Float1779Output_2287: float (5 downto -14);
Signal ProductNode_Float1780weight : float ( 5 downto -14 ) := to_float (0.780732,5,14);

Signal ProductNode_Float1780Output_2288: float (5 downto -14);
Signal ProductNode_Float1781weight : float ( 5 downto -14 ) := to_float (0.917308,5,14);

Signal ProductNode_Float1781Output_2289: float (5 downto -14);
Signal SumNode_Float508Output_2290: float (5 downto -14);
Signal ProductNode_Float1782Output_2291: float (5 downto -14);
Signal ProductNode_Float1783weight : float ( 5 downto -14 ) := to_float (0.631626,5,14);

Signal ProductNode_Float1783Output_2292: float (5 downto -14);
Signal ProductNode_Float1784weight : float ( 5 downto -14 ) := to_float (0.453222,5,14);

Signal ProductNode_Float1784Output_2293: float (5 downto -14);
Signal ProductNode_Float1785weight : float ( 5 downto -14 ) := to_float (0.996146,5,14);

Signal ProductNode_Float1785Output_2294: float (5 downto -14);
Signal SumNode_Float509Output_2295: float (5 downto -14);
Signal ProductNode_Float1786Output_2296: float (5 downto -14);
Signal ProductNode_Float1787weight : float ( 5 downto -14 ) := to_float (0.870697,5,14);

Signal ProductNode_Float1787Output_2297: float (5 downto -14);
Signal ProductNode_Float1788weight : float ( 5 downto -14 ) := to_float (0.753690,5,14);

Signal ProductNode_Float1788Output_2298: float (5 downto -14);
Signal ProductNode_Float1789weight : float ( 5 downto -14 ) := to_float (0.936763,5,14);

Signal ProductNode_Float1789Output_2299: float (5 downto -14);
Signal ProductNode_Float1790weight : float ( 5 downto -14 ) := to_float (0.870404,5,14);

Signal ProductNode_Float1790Output_2300: float (5 downto -14);
Signal ProductNode_Float1791weight : float ( 5 downto -14 ) := to_float (0.933776,5,14);

Signal ProductNode_Float1791Output_2301: float (5 downto -14);
Signal ProductNode_Float1792weight : float ( 5 downto -14 ) := to_float (0.973389,5,14);

Signal ProductNode_Float1792Output_2302: float (5 downto -14);
Signal SumNode_Float510Output_2303: float (5 downto -14);
Signal ProductNode_Float1793Output_2304: float (5 downto -14);
Signal ProductNode_Float1794weight : float ( 5 downto -14 ) := to_float (0.912549,5,14);

Signal ProductNode_Float1794Output_2305: float (5 downto -14);
Signal SumNode_Float511Output_2306: float (5 downto -14);
Signal ProductNode_Float1795Output_2307: float (5 downto -14);
Signal ProductNode_Float1796weight : float ( 5 downto -14 ) := to_float (0.658116,5,14);

Signal ProductNode_Float1796Output_2308: float (5 downto -14);
Signal ProductNode_Float1797weight : float ( 5 downto -14 ) := to_float (0.890735,5,14);

Signal ProductNode_Float1797Output_2309: float (5 downto -14);
Signal ProductNode_Float1798weight : float ( 5 downto -14 ) := to_float (0.382644,5,14);

Signal ProductNode_Float1798Output_2310: float (5 downto -14);
Signal ProductNode_Float1799weight : float ( 5 downto -14 ) := to_float (0.998354,5,14);

Signal ProductNode_Float1799Output_2311: float (5 downto -14);
Signal SumNode_Float512Output_2312: float (5 downto -14);
Signal ProductNode_Float1800Output_2313: float (5 downto -14);
Signal ProductNode_Float1801weight : float ( 5 downto -14 ) := to_float (0.551341,5,14);

Signal ProductNode_Float1801Output_2314: float (5 downto -14);
Signal ProductNode_Float1802weight : float ( 5 downto -14 ) := to_float (0.795357,5,14);

Signal ProductNode_Float1802Output_2315: float (5 downto -14);
Signal ProductNode_Float1803weight : float ( 5 downto -14 ) := to_float (0.948695,5,14);

Signal ProductNode_Float1803Output_2316: float (5 downto -14);
Signal ProductNode_Float1804weight : float ( 5 downto -14 ) := to_float (0.989597,5,14);

Signal ProductNode_Float1804Output_2317: float (5 downto -14);
Signal ProductNode_Float1805weight : float ( 5 downto -14 ) := to_float (0.577708,5,14);

Signal ProductNode_Float1805Output_2318: float (5 downto -14);
Signal ProductNode_Float1806weight : float ( 5 downto -14 ) := to_float (0.981240,5,14);

Signal ProductNode_Float1806Output_2319: float (5 downto -14);
Signal SumNode_Float513Output_2320: float (5 downto -14);
Signal ProductNode_Float1807Output_2321: float (5 downto -14);
Signal ProductNode_Float1808weight : float ( 5 downto -14 ) := to_float (0.712179,5,14);

Signal ProductNode_Float1808Output_2322: float (5 downto -14);
Signal ProductNode_Float1809weight : float ( 5 downto -14 ) := to_float (0.336149,5,14);

Signal ProductNode_Float1809Output_2323: float (5 downto -14);
Signal ProductNode_Float1810weight : float ( 5 downto -14 ) := to_float (0.999140,5,14);

Signal ProductNode_Float1810Output_2324: float (5 downto -14);
Signal SumNode_Float514Output_2325: float (5 downto -14);
Signal ProductNode_Float1811Output_2326: float (5 downto -14);
Signal ProductNode_Float1812weight : float ( 5 downto -14 ) := to_float (0.551341,5,14);

Signal ProductNode_Float1812Output_2327: float (5 downto -14);
Signal ProductNode_Float1813weight : float ( 5 downto -14 ) := to_float (0.926235,5,14);

Signal ProductNode_Float1813Output_2328: float (5 downto -14);
Signal ProductNode_Float1814weight : float ( 5 downto -14 ) := to_float (0.981519,5,14);

Signal ProductNode_Float1814Output_2329: float (5 downto -14);
Signal ProductNode_Float1815weight : float ( 5 downto -14 ) := to_float (0.989597,5,14);

Signal ProductNode_Float1815Output_2330: float (5 downto -14);
Signal ProductNode_Float1816weight : float ( 5 downto -14 ) := to_float (0.986786,5,14);

Signal ProductNode_Float1816Output_2331: float (5 downto -14);
Signal ProductNode_Float1817weight : float ( 5 downto -14 ) := to_float (0.995641,5,14);

Signal ProductNode_Float1817Output_2332: float (5 downto -14);
Signal SumNode_Float515Output_2333: float (5 downto -14);
Signal ProductNode_Float1818Output_2334: float (5 downto -14);
Signal ProductNode_Float1819weight : float ( 5 downto -14 ) := to_float (0.972670,5,14);

Signal ProductNode_Float1819Output_2335: float (5 downto -14);
Signal SumNode_Float516Output_2336: float (5 downto -14);
Signal ProductNode_Float1820Output_2337: float (5 downto -14);
Signal ProductNode_Float1821weight : float ( 5 downto -14 ) := to_float (0.531350,5,14);

Signal ProductNode_Float1821Output_2338: float (5 downto -14);
Signal SumNode_Float517Output_2339: float (5 downto -14);
Signal ProductNode_Float1822Output_2340: float (5 downto -14);
Signal ProductNode_Float1823weight : float ( 5 downto -14 ) := to_float (0.816772,5,14);

Signal ProductNode_Float1823Output_2341: float (5 downto -14);
Signal SumNode_Float518Output_2342: float (5 downto -14);
Signal ProductNode_Float1824Output_2343: float (5 downto -14);
Signal ProductNode_Float1825weight : float ( 5 downto -14 ) := to_float (0.965849,5,14);

Signal ProductNode_Float1825Output_2344: float (5 downto -14);
Signal ProductNode_Float1826weight : float ( 5 downto -14 ) := to_float (0.692695,5,14);

Signal ProductNode_Float1826Output_2345: float (5 downto -14);
Signal SumNode_Float519Output_2346: float (5 downto -14);
Signal ProductNode_Float1827Output_2347: float (5 downto -14);
Signal ProductNode_Float1828weight : float ( 5 downto -14 ) := to_float (0.880399,5,14);

Signal ProductNode_Float1828Output_2348: float (5 downto -14);
Signal ProductNode_Float1829weight : float ( 5 downto -14 ) := to_float (0.997554,5,14);

Signal ProductNode_Float1829Output_2349: float (5 downto -14);
Signal ProductNode_Float1830weight : float ( 5 downto -14 ) := to_float (0.414069,5,14);

Signal ProductNode_Float1830Output_2350: float (5 downto -14);
Signal SumNode_Float520Output_2351: float (5 downto -14);
Signal ProductNode_Float1831Output_2352: float (5 downto -14);
Signal ProductNode_Float1832weight : float ( 5 downto -14 ) := to_float (0.919660,5,14);

Signal ProductNode_Float1832Output_2353: float (5 downto -14);
Signal ProductNode_Float1833weight : float ( 5 downto -14 ) := to_float (0.806938,5,14);

Signal ProductNode_Float1833Output_2354: float (5 downto -14);
Signal SumNode_Float521Output_2355: float (5 downto -14);
Signal ProductNode_Float1834Output_2356: float (5 downto -14);
Signal ProductNode_Float1835weight : float ( 5 downto -14 ) := to_float (0.860235,5,14);

Signal ProductNode_Float1835Output_2357: float (5 downto -14);
Signal ProductNode_Float1836weight : float ( 5 downto -14 ) := to_float (0.989739,5,14);

Signal ProductNode_Float1836Output_2358: float (5 downto -14);
Signal ProductNode_Float1837weight : float ( 5 downto -14 ) := to_float (0.549861,5,14);

Signal ProductNode_Float1837Output_2359: float (5 downto -14);
Signal SumNode_Float522Output_2360: float (5 downto -14);
Signal ProductNode_Float1838Output_2361: float (5 downto -14);
Signal SumNode_Float523Output_2362: float (5 downto -14);
Signal ProductNode_Float1839Output_2363: float (5 downto -14);
Signal ProductNode_Float1840weight : float ( 5 downto -14 ) := to_float (0.984104,5,14);

Signal ProductNode_Float1840Output_2364: float (5 downto -14);
Signal ProductNode_Float1841weight : float ( 5 downto -14 ) := to_float (0.793165,5,14);

Signal ProductNode_Float1841Output_2365: float (5 downto -14);
Signal ProductNode_Float1842weight : float ( 5 downto -14 ) := to_float (0.927417,5,14);

Signal ProductNode_Float1842Output_2366: float (5 downto -14);
Signal SumNode_Float524Output_2367: float (5 downto -14);
Signal ProductNode_Float1843Output_2368: float (5 downto -14);
Signal ProductNode_Float1844weight : float ( 5 downto -14 ) := to_float (0.726095,5,14);

Signal ProductNode_Float1844Output_2369: float (5 downto -14);
Signal ProductNode_Float1845weight : float ( 5 downto -14 ) := to_float (0.988880,5,14);

Signal ProductNode_Float1845Output_2370: float (5 downto -14);
Signal ProductNode_Float1846weight : float ( 5 downto -14 ) := to_float (0.558577,5,14);

Signal ProductNode_Float1846Output_2371: float (5 downto -14);
Signal SumNode_Float525Output_2372: float (5 downto -14);
Signal ProductNode_Float1847Output_2373: float (5 downto -14);
Signal ProductNode_Float1848weight : float ( 5 downto -14 ) := to_float (0.649155,5,14);

Signal ProductNode_Float1848Output_2374: float (5 downto -14);
Signal ProductNode_Float1849weight : float ( 5 downto -14 ) := to_float (0.975801,5,14);

Signal ProductNode_Float1849Output_2375: float (5 downto -14);
Signal SumNode_Float526Output_2376: float (5 downto -14);
Signal ProductNode_Float1850Output_2377: float (5 downto -14);
Signal ProductNode_Float1851weight : float ( 5 downto -14 ) := to_float (0.955917,5,14);

Signal ProductNode_Float1851Output_2378: float (5 downto -14);
Signal ProductNode_Float1852weight : float ( 5 downto -14 ) := to_float (0.985013,5,14);

Signal ProductNode_Float1852Output_2379: float (5 downto -14);
Signal ProductNode_Float1853weight : float ( 5 downto -14 ) := to_float (0.592017,5,14);

Signal ProductNode_Float1853Output_2380: float (5 downto -14);
Signal SumNode_Float527Output_2381: float (5 downto -14);
Signal ProductNode_Float1854Output_2382: float (5 downto -14);
Signal SumNode_Float528Output_2383: float (5 downto -14);
Signal ProductNode_Float1855Output_2384: float (5 downto -14);
Signal ProductNode_Float1856weight : float ( 5 downto -14 ) := to_float (0.598812,5,14);

Signal ProductNode_Float1856Output_2385: float (5 downto -14);
Signal SumNode_Float529Output_2386: float (5 downto -14);
Signal ProductNode_Float1857Output_2387: float (5 downto -14);
Signal ProductNode_Float1858weight : float ( 5 downto -14 ) := to_float (0.807423,5,14);

Signal ProductNode_Float1858Output_2388: float (5 downto -14);
Signal ProductNode_Float1859weight : float ( 5 downto -14 ) := to_float (0.919372,5,14);

Signal ProductNode_Float1859Output_2389: float (5 downto -14);
Signal SumNode_Float530Output_2390: float (5 downto -14);
Signal ProductNode_Float1860Output_2391: float (5 downto -14);
Signal ProductNode_Float1861weight : float ( 5 downto -14 ) := to_float (0.694473,5,14);

Signal ProductNode_Float1861Output_2392: float (5 downto -14);
Signal ProductNode_Float1862weight : float ( 5 downto -14 ) := to_float (0.843444,5,14);

Signal ProductNode_Float1862Output_2393: float (5 downto -14);
Signal ProductNode_Float1863weight : float ( 5 downto -14 ) := to_float (0.682797,5,14);

Signal ProductNode_Float1863Output_2394: float (5 downto -14);
Signal ProductNode_Float1864weight : float ( 5 downto -14 ) := to_float (0.968381,5,14);

Signal ProductNode_Float1864Output_2395: float (5 downto -14);
Signal SumNode_Float531Output_2396: float (5 downto -14);
Signal ProductNode_Float1865Output_2397: float (5 downto -14);
Signal ProductNode_Float1866weight : float ( 5 downto -14 ) := to_float (0.965376,5,14);

Signal ProductNode_Float1866Output_2398: float (5 downto -14);
Signal ProductNode_Float1867weight : float ( 5 downto -14 ) := to_float (0.697447,5,14);

Signal ProductNode_Float1867Output_2399: float (5 downto -14);
Signal SumNode_Float532Output_2400: float (5 downto -14);
Signal ProductNode_Float1868Output_2401: float (5 downto -14);
Signal ProductNode_Float1869weight : float ( 5 downto -14 ) := to_float (0.965849,5,14);

Signal ProductNode_Float1869Output_2402: float (5 downto -14);
Signal ProductNode_Float1870weight : float ( 5 downto -14 ) := to_float (0.692695,5,14);

Signal ProductNode_Float1870Output_2403: float (5 downto -14);
Signal SumNode_Float533Output_2404: float (5 downto -14);
Signal ProductNode_Float1871Output_2405: float (5 downto -14);
Signal ProductNode_Float1872weight : float ( 5 downto -14 ) := to_float (0.880399,5,14);

Signal ProductNode_Float1872Output_2406: float (5 downto -14);
Signal ProductNode_Float1873weight : float ( 5 downto -14 ) := to_float (0.997554,5,14);

Signal ProductNode_Float1873Output_2407: float (5 downto -14);
Signal ProductNode_Float1874weight : float ( 5 downto -14 ) := to_float (0.414069,5,14);

Signal ProductNode_Float1874Output_2408: float (5 downto -14);
Signal SumNode_Float534Output_2409: float (5 downto -14);
Signal ProductNode_Float1875Output_2410: float (5 downto -14);
Signal ProductNode_Float1876weight : float ( 5 downto -14 ) := to_float (0.919660,5,14);

Signal ProductNode_Float1876Output_2411: float (5 downto -14);
Signal ProductNode_Float1877weight : float ( 5 downto -14 ) := to_float (0.806938,5,14);

Signal ProductNode_Float1877Output_2412: float (5 downto -14);
Signal SumNode_Float535Output_2413: float (5 downto -14);
Signal ProductNode_Float1878Output_2414: float (5 downto -14);
Signal ProductNode_Float1879weight : float ( 5 downto -14 ) := to_float (0.860235,5,14);

Signal ProductNode_Float1879Output_2415: float (5 downto -14);
Signal ProductNode_Float1880weight : float ( 5 downto -14 ) := to_float (0.989739,5,14);

Signal ProductNode_Float1880Output_2416: float (5 downto -14);
Signal ProductNode_Float1881weight : float ( 5 downto -14 ) := to_float (0.549861,5,14);

Signal ProductNode_Float1881Output_2417: float (5 downto -14);
Signal SumNode_Float536Output_2418: float (5 downto -14);
Signal ProductNode_Float1882Output_2419: float (5 downto -14);
Signal SumNode_Float537Output_2420: float (5 downto -14);
Signal ProductNode_Float1883Output_2421: float (5 downto -14);
Signal ProductNode_Float1884weight : float ( 5 downto -14 ) := to_float (0.932937,5,14);

Signal ProductNode_Float1884Output_2422: float (5 downto -14);
Signal ProductNode_Float1885weight : float ( 5 downto -14 ) := to_float (0.793165,5,14);

Signal ProductNode_Float1885Output_2423: float (5 downto -14);
Signal ProductNode_Float1886weight : float ( 5 downto -14 ) := to_float (0.927417,5,14);

Signal ProductNode_Float1886Output_2424: float (5 downto -14);
Signal SumNode_Float538Output_2425: float (5 downto -14);
Signal ProductNode_Float1887Output_2426: float (5 downto -14);
Signal ProductNode_Float1888weight : float ( 5 downto -14 ) := to_float (0.726095,5,14);

Signal ProductNode_Float1888Output_2427: float (5 downto -14);
Signal ProductNode_Float1889weight : float ( 5 downto -14 ) := to_float (0.988880,5,14);

Signal ProductNode_Float1889Output_2428: float (5 downto -14);
Signal ProductNode_Float1890weight : float ( 5 downto -14 ) := to_float (0.558577,5,14);

Signal ProductNode_Float1890Output_2429: float (5 downto -14);
Signal SumNode_Float539Output_2430: float (5 downto -14);
Signal ProductNode_Float1891Output_2431: float (5 downto -14);
Signal ProductNode_Float1892weight : float ( 5 downto -14 ) := to_float (0.649155,5,14);

Signal ProductNode_Float1892Output_2432: float (5 downto -14);
Signal ProductNode_Float1893weight : float ( 5 downto -14 ) := to_float (0.975801,5,14);

Signal ProductNode_Float1893Output_2433: float (5 downto -14);
Signal SumNode_Float540Output_2434: float (5 downto -14);
Signal ProductNode_Float1894Output_2435: float (5 downto -14);
Signal ProductNode_Float1895weight : float ( 5 downto -14 ) := to_float (0.955917,5,14);

Signal ProductNode_Float1895Output_2436: float (5 downto -14);
Signal ProductNode_Float1896weight : float ( 5 downto -14 ) := to_float (0.985013,5,14);

Signal ProductNode_Float1896Output_2437: float (5 downto -14);
Signal ProductNode_Float1897weight : float ( 5 downto -14 ) := to_float (0.592017,5,14);

Signal ProductNode_Float1897Output_2438: float (5 downto -14);
Signal SumNode_Float541Output_2439: float (5 downto -14);
Signal ProductNode_Float1898Output_2440: float (5 downto -14);
Signal SumNode_Float542Output_2441: float (5 downto -14);
Signal ProductNode_Float1899Output_2442: float (5 downto -14);
Signal ProductNode_Float1900weight : float ( 5 downto -14 ) := to_float (0.782438,5,14);

Signal ProductNode_Float1900Output_2443: float (5 downto -14);
Signal SumNode_Float543Output_2444: float (5 downto -14);
Signal ProductNode_Float1901Output_2445: float (5 downto -14);
Signal ProductNode_Float1902weight : float ( 5 downto -14 ) := to_float (0.623360,5,14);

Signal ProductNode_Float1902Output_2446: float (5 downto -14);
Signal ProductNode_Float1903weight : float ( 5 downto -14 ) := to_float (0.980424,5,14);

Signal ProductNode_Float1903Output_2447: float (5 downto -14);
Signal SumNode_Float544Output_2448: float (5 downto -14);
Signal ProductNode_Float1904Output_2449: float (5 downto -14);
Signal ProductNode_Float1905weight : float ( 5 downto -14 ) := to_float (0.694473,5,14);

Signal ProductNode_Float1905Output_2450: float (5 downto -14);
Signal ProductNode_Float1906weight : float ( 5 downto -14 ) := to_float (0.894649,5,14);

Signal ProductNode_Float1906Output_2451: float (5 downto -14);
Signal ProductNode_Float1907weight : float ( 5 downto -14 ) := to_float (0.482891,5,14);

Signal ProductNode_Float1907Output_2452: float (5 downto -14);
Signal ProductNode_Float1908weight : float ( 5 downto -14 ) := to_float (0.994693,5,14);

Signal ProductNode_Float1908Output_2453: float (5 downto -14);
Signal SumNode_Float545Output_2454: float (5 downto -14);
Signal ProductNode_Float1909Output_2455: float (5 downto -14);
Signal ProductNode_Float1910weight : float ( 5 downto -14 ) := to_float (0.965376,5,14);

Signal ProductNode_Float1910Output_2456: float (5 downto -14);
Signal ProductNode_Float1911weight : float ( 5 downto -14 ) := to_float (0.964572,5,14);

Signal ProductNode_Float1911Output_2457: float (5 downto -14);
Signal SumNode_Float546Output_2458: float (5 downto -14);
Signal ProductNode_Float1912Output_2459: float (5 downto -14);
Signal SumNode_Float547Output_2460: float (5 downto -14);
Signal ProductNode_Float1913Output_2461: float (5 downto -14);
Signal ProductNode_Float1914weight : float ( 5 downto -14 ) := to_float (0.926565,5,14);

Signal ProductNode_Float1914Output_2462: float (5 downto -14);
Signal ProductNode_Float1915weight : float ( 5 downto -14 ) := to_float (0.965849,5,14);

Signal ProductNode_Float1915Output_2463: float (5 downto -14);
Signal ProductNode_Float1916weight : float ( 5 downto -14 ) := to_float (0.692695,5,14);

Signal ProductNode_Float1916Output_2464: float (5 downto -14);
Signal SumNode_Float548Output_2465: float (5 downto -14);
Signal ProductNode_Float1917Output_2466: float (5 downto -14);
Signal ProductNode_Float1918weight : float ( 5 downto -14 ) := to_float (0.880399,5,14);

Signal ProductNode_Float1918Output_2467: float (5 downto -14);
Signal ProductNode_Float1919weight : float ( 5 downto -14 ) := to_float (0.966381,5,14);

Signal ProductNode_Float1919Output_2468: float (5 downto -14);
Signal ProductNode_Float1920weight : float ( 5 downto -14 ) := to_float (0.690672,5,14);

Signal ProductNode_Float1920Output_2469: float (5 downto -14);
Signal SumNode_Float549Output_2470: float (5 downto -14);
Signal ProductNode_Float1921Output_2471: float (5 downto -14);
Signal ProductNode_Float1922weight : float ( 5 downto -14 ) := to_float (0.919660,5,14);

Signal ProductNode_Float1922Output_2472: float (5 downto -14);
Signal ProductNode_Float1923weight : float ( 5 downto -14 ) := to_float (0.806938,5,14);

Signal ProductNode_Float1923Output_2473: float (5 downto -14);
Signal SumNode_Float550Output_2474: float (5 downto -14);
Signal ProductNode_Float1924Output_2475: float (5 downto -14);
Signal ProductNode_Float1925weight : float ( 5 downto -14 ) := to_float (0.860235,5,14);

Signal ProductNode_Float1925Output_2476: float (5 downto -14);
Signal ProductNode_Float1926weight : float ( 5 downto -14 ) := to_float (0.941870,5,14);

Signal ProductNode_Float1926Output_2477: float (5 downto -14);
Signal ProductNode_Float1927weight : float ( 5 downto -14 ) := to_float (0.763101,5,14);

Signal ProductNode_Float1927Output_2478: float (5 downto -14);
Signal SumNode_Float551Output_2479: float (5 downto -14);
Signal ProductNode_Float1928Output_2480: float (5 downto -14);
Signal SumNode_Float552Output_2481: float (5 downto -14);
Signal ProductNode_Float1929Output_2482: float (5 downto -14);
Signal ProductNode_Float1930weight : float ( 5 downto -14 ) := to_float (0.924413,5,14);

Signal ProductNode_Float1930Output_2483: float (5 downto -14);
Signal ProductNode_Float1931weight : float ( 5 downto -14 ) := to_float (0.793165,5,14);

Signal ProductNode_Float1931Output_2484: float (5 downto -14);
Signal ProductNode_Float1932weight : float ( 5 downto -14 ) := to_float (0.927417,5,14);

Signal ProductNode_Float1932Output_2485: float (5 downto -14);
Signal SumNode_Float553Output_2486: float (5 downto -14);
Signal ProductNode_Float1933Output_2487: float (5 downto -14);
Signal ProductNode_Float1934weight : float ( 5 downto -14 ) := to_float (0.726095,5,14);

Signal ProductNode_Float1934Output_2488: float (5 downto -14);
Signal ProductNode_Float1935weight : float ( 5 downto -14 ) := to_float (0.909585,5,14);

Signal ProductNode_Float1935Output_2489: float (5 downto -14);
Signal ProductNode_Float1936weight : float ( 5 downto -14 ) := to_float (0.822920,5,14);

Signal ProductNode_Float1936Output_2490: float (5 downto -14);
Signal SumNode_Float554Output_2491: float (5 downto -14);
Signal ProductNode_Float1937Output_2492: float (5 downto -14);
Signal ProductNode_Float1938weight : float ( 5 downto -14 ) := to_float (0.649155,5,14);

Signal ProductNode_Float1938Output_2493: float (5 downto -14);
Signal ProductNode_Float1939weight : float ( 5 downto -14 ) := to_float (0.975801,5,14);

Signal ProductNode_Float1939Output_2494: float (5 downto -14);
Signal SumNode_Float555Output_2495: float (5 downto -14);
Signal ProductNode_Float1940Output_2496: float (5 downto -14);
Signal ProductNode_Float1941weight : float ( 5 downto -14 ) := to_float (0.955917,5,14);

Signal ProductNode_Float1941Output_2497: float (5 downto -14);
Signal ProductNode_Float1942weight : float ( 5 downto -14 ) := to_float (0.790147,5,14);

Signal ProductNode_Float1942Output_2498: float (5 downto -14);
Signal ProductNode_Float1943weight : float ( 5 downto -14 ) := to_float (0.929014,5,14);

Signal ProductNode_Float1943Output_2499: float (5 downto -14);
Signal SumNode_Float556Output_2500: float (5 downto -14);
Signal ProductNode_Float1944Output_2501: float (5 downto -14);
Signal SumNode_Float557Output_2502: float (5 downto -14);
Signal ProductNode_Float1945Output_2503: float (5 downto -14);
Signal ProductNode_Float1946weight : float ( 5 downto -14 ) := to_float (0.798666,5,14);

Signal ProductNode_Float1946Output_2504: float (5 downto -14);
Signal SumNode_Float558Output_2505: float (5 downto -14);
Signal ProductNode_Float1947Output_2506: float (5 downto -14);
Signal ProductNode_Float1948weight : float ( 5 downto -14 ) := to_float (0.807423,5,14);

Signal ProductNode_Float1948Output_2507: float (5 downto -14);
Signal ProductNode_Float1949weight : float ( 5 downto -14 ) := to_float (0.919372,5,14);

Signal ProductNode_Float1949Output_2508: float (5 downto -14);
Signal SumNode_Float559Output_2509: float (5 downto -14);
Signal ProductNode_Float1950Output_2510: float (5 downto -14);
Signal ProductNode_Float1951weight : float ( 5 downto -14 ) := to_float (0.579487,5,14);

Signal ProductNode_Float1951Output_2511: float (5 downto -14);
Signal ProductNode_Float1952weight : float ( 5 downto -14 ) := to_float (0.790558,5,14);

Signal ProductNode_Float1952Output_2512: float (5 downto -14);
Signal ProductNode_Float1953weight : float ( 5 downto -14 ) := to_float (0.682797,5,14);

Signal ProductNode_Float1953Output_2513: float (5 downto -14);
Signal ProductNode_Float1954weight : float ( 5 downto -14 ) := to_float (0.968381,5,14);

Signal ProductNode_Float1954Output_2514: float (5 downto -14);
Signal SumNode_Float560Output_2515: float (5 downto -14);
Signal ProductNode_Float1955Output_2516: float (5 downto -14);
Signal ProductNode_Float1956weight : float ( 5 downto -14 ) := to_float (0.986575,5,14);

Signal ProductNode_Float1956Output_2517: float (5 downto -14);
Signal ProductNode_Float1957weight : float ( 5 downto -14 ) := to_float (0.578242,5,14);

Signal ProductNode_Float1957Output_2518: float (5 downto -14);
Signal SumNode_Float561Output_2519: float (5 downto -14);
Signal ProductNode_Float1958Output_2520: float (5 downto -14);
Signal ProductNode_Float1959weight : float ( 5 downto -14 ) := to_float (0.965849,5,14);

Signal ProductNode_Float1959Output_2521: float (5 downto -14);
Signal ProductNode_Float1960weight : float ( 5 downto -14 ) := to_float (0.692695,5,14);

Signal ProductNode_Float1960Output_2522: float (5 downto -14);
Signal SumNode_Float562Output_2523: float (5 downto -14);
Signal ProductNode_Float1961Output_2524: float (5 downto -14);
Signal ProductNode_Float1962weight : float ( 5 downto -14 ) := to_float (0.880399,5,14);

Signal ProductNode_Float1962Output_2525: float (5 downto -14);
Signal ProductNode_Float1963weight : float ( 5 downto -14 ) := to_float (0.966381,5,14);

Signal ProductNode_Float1963Output_2526: float (5 downto -14);
Signal ProductNode_Float1964weight : float ( 5 downto -14 ) := to_float (0.690672,5,14);

Signal ProductNode_Float1964Output_2527: float (5 downto -14);
Signal SumNode_Float563Output_2528: float (5 downto -14);
Signal ProductNode_Float1965Output_2529: float (5 downto -14);
Signal ProductNode_Float1966weight : float ( 5 downto -14 ) := to_float (0.919660,5,14);

Signal ProductNode_Float1966Output_2530: float (5 downto -14);
Signal ProductNode_Float1967weight : float ( 5 downto -14 ) := to_float (0.806938,5,14);

Signal ProductNode_Float1967Output_2531: float (5 downto -14);
Signal SumNode_Float564Output_2532: float (5 downto -14);
Signal ProductNode_Float1968Output_2533: float (5 downto -14);
Signal ProductNode_Float1969weight : float ( 5 downto -14 ) := to_float (0.860235,5,14);

Signal ProductNode_Float1969Output_2534: float (5 downto -14);
Signal ProductNode_Float1970weight : float ( 5 downto -14 ) := to_float (0.941870,5,14);

Signal ProductNode_Float1970Output_2535: float (5 downto -14);
Signal ProductNode_Float1971weight : float ( 5 downto -14 ) := to_float (0.763101,5,14);

Signal ProductNode_Float1971Output_2536: float (5 downto -14);
Signal SumNode_Float565Output_2537: float (5 downto -14);
Signal ProductNode_Float1972Output_2538: float (5 downto -14);
Signal SumNode_Float566Output_2539: float (5 downto -14);
Signal ProductNode_Float1973Output_2540: float (5 downto -14);
Signal ProductNode_Float1974weight : float ( 5 downto -14 ) := to_float (0.693688,5,14);

Signal ProductNode_Float1974Output_2541: float (5 downto -14);
Signal ProductNode_Float1975weight : float ( 5 downto -14 ) := to_float (0.793165,5,14);

Signal ProductNode_Float1975Output_2542: float (5 downto -14);
Signal ProductNode_Float1976weight : float ( 5 downto -14 ) := to_float (0.927417,5,14);

Signal ProductNode_Float1976Output_2543: float (5 downto -14);
Signal SumNode_Float567Output_2544: float (5 downto -14);
Signal ProductNode_Float1977Output_2545: float (5 downto -14);
Signal ProductNode_Float1978weight : float ( 5 downto -14 ) := to_float (0.726095,5,14);

Signal ProductNode_Float1978Output_2546: float (5 downto -14);
Signal ProductNode_Float1979weight : float ( 5 downto -14 ) := to_float (0.909585,5,14);

Signal ProductNode_Float1979Output_2547: float (5 downto -14);
Signal ProductNode_Float1980weight : float ( 5 downto -14 ) := to_float (0.822920,5,14);

Signal ProductNode_Float1980Output_2548: float (5 downto -14);
Signal SumNode_Float568Output_2549: float (5 downto -14);
Signal ProductNode_Float1981Output_2550: float (5 downto -14);
Signal ProductNode_Float1982weight : float ( 5 downto -14 ) := to_float (0.649155,5,14);

Signal ProductNode_Float1982Output_2551: float (5 downto -14);
Signal ProductNode_Float1983weight : float ( 5 downto -14 ) := to_float (0.975801,5,14);

Signal ProductNode_Float1983Output_2552: float (5 downto -14);
Signal SumNode_Float569Output_2553: float (5 downto -14);
Signal ProductNode_Float1984Output_2554: float (5 downto -14);
Signal ProductNode_Float1985weight : float ( 5 downto -14 ) := to_float (0.955917,5,14);

Signal ProductNode_Float1985Output_2555: float (5 downto -14);
Signal ProductNode_Float1986weight : float ( 5 downto -14 ) := to_float (0.790147,5,14);

Signal ProductNode_Float1986Output_2556: float (5 downto -14);
Signal ProductNode_Float1987weight : float ( 5 downto -14 ) := to_float (0.929014,5,14);

Signal ProductNode_Float1987Output_2557: float (5 downto -14);
Signal SumNode_Float570Output_2558: float (5 downto -14);
Signal ProductNode_Float1988Output_2559: float (5 downto -14);
Signal SumNode_Float571Output_2560: float (5 downto -14);
Signal ProductNode_Float1989Output_2561: float (5 downto -14);
Signal ProductNode_Float1990weight : float ( 5 downto -14 ) := to_float (0.965586,5,14);

Signal ProductNode_Float1990Output_2562: float (5 downto -14);
Signal SumNode_Float572Output_2563: float (5 downto -14);
Signal ProductNode_Float1991Output_2564: float (5 downto -14);
Signal ProductNode_Float1992weight : float ( 5 downto -14 ) := to_float (0.623360,5,14);

Signal ProductNode_Float1992Output_2565: float (5 downto -14);
Signal ProductNode_Float1993weight : float ( 5 downto -14 ) := to_float (0.980424,5,14);

Signal ProductNode_Float1993Output_2566: float (5 downto -14);
Signal SumNode_Float573Output_2567: float (5 downto -14);
Signal ProductNode_Float1994Output_2568: float (5 downto -14);
Signal ProductNode_Float1995weight : float ( 5 downto -14 ) := to_float (0.579487,5,14);

Signal ProductNode_Float1995Output_2569: float (5 downto -14);
Signal ProductNode_Float1996weight : float ( 5 downto -14 ) := to_float (0.928799,5,14);

Signal ProductNode_Float1996Output_2570: float (5 downto -14);
Signal ProductNode_Float1997weight : float ( 5 downto -14 ) := to_float (0.482891,5,14);

Signal ProductNode_Float1997Output_2571: float (5 downto -14);
Signal ProductNode_Float1998weight : float ( 5 downto -14 ) := to_float (0.994693,5,14);

Signal ProductNode_Float1998Output_2572: float (5 downto -14);
Signal SumNode_Float574Output_2573: float (5 downto -14);
Signal ProductNode_Float1999Output_2574: float (5 downto -14);
Signal ProductNode_Float2000weight : float ( 5 downto -14 ) := to_float (0.986575,5,14);

Signal ProductNode_Float2000Output_2575: float (5 downto -14);
Signal ProductNode_Float2001weight : float ( 5 downto -14 ) := to_float (0.986723,5,14);

Signal ProductNode_Float2001Output_2576: float (5 downto -14);
Signal SumNode_Float575Output_2577: float (5 downto -14);
Signal ProductNode_Float2002Output_2578: float (5 downto -14);
Signal SumNode_Float576Output_2579: float (5 downto -14);
Signal ProductNode_Float2003Output_2580: float (5 downto -14);
Signal ProductNode_Float2004weight : float ( 5 downto -14 ) := to_float (0.794749,5,14);

Signal ProductNode_Float2004Output_2581: float (5 downto -14);
Signal SumNode_Float577Output_2582: float (5 downto -14);
Signal ProductNode_Float2005Output_2583: float (5 downto -14);
Signal ProductNode_Float2006weight : float ( 5 downto -14 ) := to_float (0.848299,5,14);

Signal ProductNode_Float2006Output_2584: float (5 downto -14);
Signal ProductNode_Float2007weight : float ( 5 downto -14 ) := to_float (0.895308,5,14);

Signal ProductNode_Float2007Output_2585: float (5 downto -14);
Signal ProductNode_Float2008weight : float ( 5 downto -14 ) := to_float (0.842608,5,14);

Signal ProductNode_Float2008Output_2586: float (5 downto -14);
Signal SumNode_Float578Output_2587: float (5 downto -14);
Signal ProductNode_Float2009Output_2588: float (5 downto -14);
Signal ProductNode_Float2010weight : float ( 5 downto -14 ) := to_float (0.870697,5,14);

Signal ProductNode_Float2010Output_2589: float (5 downto -14);
Signal ProductNode_Float2011weight : float ( 5 downto -14 ) := to_float (0.945793,5,14);

Signal ProductNode_Float2011Output_2590: float (5 downto -14);
Signal ProductNode_Float2012weight : float ( 5 downto -14 ) := to_float (0.954870,5,14);

Signal ProductNode_Float2012Output_2591: float (5 downto -14);
Signal ProductNode_Float2013weight : float ( 5 downto -14 ) := to_float (0.870404,5,14);

Signal ProductNode_Float2013Output_2592: float (5 downto -14);
Signal ProductNode_Float2014weight : float ( 5 downto -14 ) := to_float (0.780732,5,14);

Signal ProductNode_Float2014Output_2593: float (5 downto -14);
Signal ProductNode_Float2015weight : float ( 5 downto -14 ) := to_float (0.810846,5,14);

Signal ProductNode_Float2015Output_2594: float (5 downto -14);
Signal SumNode_Float579Output_2595: float (5 downto -14);
Signal ProductNode_Float2016Output_2596: float (5 downto -14);
Signal ProductNode_Float2017weight : float ( 5 downto -14 ) := to_float (0.531606,5,14);

Signal ProductNode_Float2017Output_2597: float (5 downto -14);
Signal ProductNode_Float2018weight : float ( 5 downto -14 ) := to_float (0.669241,5,14);

Signal ProductNode_Float2018Output_2598: float (5 downto -14);
Signal ProductNode_Float2019weight : float ( 5 downto -14 ) := to_float (0.971580,5,14);

Signal ProductNode_Float2019Output_2599: float (5 downto -14);
Signal SumNode_Float580Output_2600: float (5 downto -14);
Signal ProductNode_Float2020Output_2601: float (5 downto -14);
Signal ProductNode_Float2021weight : float ( 5 downto -14 ) := to_float (0.870697,5,14);

Signal ProductNode_Float2021Output_2602: float (5 downto -14);
Signal ProductNode_Float2022weight : float ( 5 downto -14 ) := to_float (0.753690,5,14);

Signal ProductNode_Float2022Output_2603: float (5 downto -14);
Signal ProductNode_Float2023weight : float ( 5 downto -14 ) := to_float (0.774480,5,14);

Signal ProductNode_Float2023Output_2604: float (5 downto -14);
Signal ProductNode_Float2024weight : float ( 5 downto -14 ) := to_float (0.870404,5,14);

Signal ProductNode_Float2024Output_2605: float (5 downto -14);
Signal ProductNode_Float2025weight : float ( 5 downto -14 ) := to_float (0.933776,5,14);

Signal ProductNode_Float2025Output_2606: float (5 downto -14);
Signal ProductNode_Float2026weight : float ( 5 downto -14 ) := to_float (0.660973,5,14);

Signal ProductNode_Float2026Output_2607: float (5 downto -14);
Signal SumNode_Float581Output_2608: float (5 downto -14);
Signal ProductNode_Float2027Output_2609: float (5 downto -14);
Signal ProductNode_Float2028weight : float ( 5 downto -14 ) := to_float (0.870862,5,14);

Signal ProductNode_Float2028Output_2610: float (5 downto -14);
Signal SumNode_Float582Output_2611: float (5 downto -14);
Signal ProductNode_Float2029Output_2612: float (5 downto -14);
Signal ProductNode_Float2030weight : float ( 5 downto -14 ) := to_float (0.888715,5,14);

Signal ProductNode_Float2030Output_2613: float (5 downto -14);
Signal ProductNode_Float2031weight : float ( 5 downto -14 ) := to_float (0.890735,5,14);

Signal ProductNode_Float2031Output_2614: float (5 downto -14);
Signal ProductNode_Float2032weight : float ( 5 downto -14 ) := to_float (0.689002,5,14);

Signal ProductNode_Float2032Output_2615: float (5 downto -14);
Signal ProductNode_Float2033weight : float ( 5 downto -14 ) := to_float (0.966814,5,14);

Signal ProductNode_Float2033Output_2616: float (5 downto -14);
Signal SumNode_Float583Output_2617: float (5 downto -14);
Signal ProductNode_Float2034Output_2618: float (5 downto -14);
Signal ProductNode_Float2035weight : float ( 5 downto -14 ) := to_float (0.551341,5,14);

Signal ProductNode_Float2035Output_2619: float (5 downto -14);
Signal ProductNode_Float2036weight : float ( 5 downto -14 ) := to_float (0.795357,5,14);

Signal ProductNode_Float2036Output_2620: float (5 downto -14);
Signal ProductNode_Float2037weight : float ( 5 downto -14 ) := to_float (0.746308,5,14);

Signal ProductNode_Float2037Output_2621: float (5 downto -14);
Signal ProductNode_Float2038weight : float ( 5 downto -14 ) := to_float (0.989597,5,14);

Signal ProductNode_Float2038Output_2622: float (5 downto -14);
Signal ProductNode_Float2039weight : float ( 5 downto -14 ) := to_float (0.577708,5,14);

Signal ProductNode_Float2039Output_2623: float (5 downto -14);
Signal ProductNode_Float2040weight : float ( 5 downto -14 ) := to_float (0.618274,5,14);

Signal ProductNode_Float2040Output_2624: float (5 downto -14);
Signal SumNode_Float584Output_2625: float (5 downto -14);
Signal ProductNode_Float2041Output_2626: float (5 downto -14);
Signal ProductNode_Float2042weight : float ( 5 downto -14 ) := to_float (0.735141,5,14);

Signal ProductNode_Float2042Output_2627: float (5 downto -14);
Signal ProductNode_Float2043weight : float ( 5 downto -14 ) := to_float (0.495915,5,14);

Signal ProductNode_Float2043Output_2628: float (5 downto -14);
Signal ProductNode_Float2044weight : float ( 5 downto -14 ) := to_float (0.993928,5,14);

Signal ProductNode_Float2044Output_2629: float (5 downto -14);
Signal SumNode_Float585Output_2630: float (5 downto -14);
Signal ProductNode_Float2045Output_2631: float (5 downto -14);
Signal ProductNode_Float2046weight : float ( 5 downto -14 ) := to_float (0.551341,5,14);

Signal ProductNode_Float2046Output_2632: float (5 downto -14);
Signal ProductNode_Float2047weight : float ( 5 downto -14 ) := to_float (0.926235,5,14);

Signal ProductNode_Float2047Output_2633: float (5 downto -14);
Signal ProductNode_Float2048weight : float ( 5 downto -14 ) := to_float (0.616494,5,14);

Signal ProductNode_Float2048Output_2634: float (5 downto -14);
Signal ProductNode_Float2049weight : float ( 5 downto -14 ) := to_float (0.989597,5,14);

Signal ProductNode_Float2049Output_2635: float (5 downto -14);
Signal ProductNode_Float2050weight : float ( 5 downto -14 ) := to_float (0.986786,5,14);

Signal ProductNode_Float2050Output_2636: float (5 downto -14);
Signal ProductNode_Float2051weight : float ( 5 downto -14 ) := to_float (0.464416,5,14);

Signal ProductNode_Float2051Output_2637: float (5 downto -14);
Signal SumNode_Float586Output_2638: float (5 downto -14);
Signal ProductNode_Float2052Output_2639: float (5 downto -14);
Signal ProductNode_Float2053weight : float ( 5 downto -14 ) := to_float (0.938375,5,14);

Signal ProductNode_Float2053Output_2640: float (5 downto -14);
Signal SumNode_Float587Output_2641: float (5 downto -14);
Signal ProductNode_Float2054Output_2642: float (5 downto -14);
Signal ProductNode_Float2055weight : float ( 5 downto -14 ) := to_float (0.978422,5,14);

Signal ProductNode_Float2055Output_2643: float (5 downto -14);
Signal SumNode_Float588Output_2644: float (5 downto -14);
Signal ProductNode_Float2056Output_2645: float (5 downto -14);
Signal ProductNode_Float2057weight : float ( 5 downto -14 ) := to_float (0.937366,5,14);

Signal ProductNode_Float2057Output_2646: float (5 downto -14);
Signal ProductNode_Float2058weight : float ( 5 downto -14 ) := to_float (0.848299,5,14);

Signal ProductNode_Float2058Output_2647: float (5 downto -14);
Signal ProductNode_Float2059weight : float ( 5 downto -14 ) := to_float (0.562709,5,14);

Signal ProductNode_Float2059Output_2648: float (5 downto -14);
Signal ProductNode_Float2060weight : float ( 5 downto -14 ) := to_float (0.988453,5,14);

Signal ProductNode_Float2060Output_2649: float (5 downto -14);
Signal SumNode_Float589Output_2650: float (5 downto -14);
Signal ProductNode_Float2061Output_2651: float (5 downto -14);
Signal ProductNode_Float2062weight : float ( 5 downto -14 ) := to_float (0.870697,5,14);

Signal ProductNode_Float2062Output_2652: float (5 downto -14);
Signal ProductNode_Float2063weight : float ( 5 downto -14 ) := to_float (0.945793,5,14);

Signal ProductNode_Float2063Output_2653: float (5 downto -14);
Signal ProductNode_Float2064weight : float ( 5 downto -14 ) := to_float (0.729204,5,14);

Signal ProductNode_Float2064Output_2654: float (5 downto -14);
Signal ProductNode_Float2065weight : float ( 5 downto -14 ) := to_float (0.870404,5,14);

Signal ProductNode_Float2065Output_2655: float (5 downto -14);
Signal ProductNode_Float2066weight : float ( 5 downto -14 ) := to_float (0.780732,5,14);

Signal ProductNode_Float2066Output_2656: float (5 downto -14);
Signal ProductNode_Float2067weight : float ( 5 downto -14 ) := to_float (0.917308,5,14);

Signal ProductNode_Float2067Output_2657: float (5 downto -14);
Signal SumNode_Float590Output_2658: float (5 downto -14);
Signal ProductNode_Float2068Output_2659: float (5 downto -14);
Signal ProductNode_Float2069weight : float ( 5 downto -14 ) := to_float (0.631626,5,14);

Signal ProductNode_Float2069Output_2660: float (5 downto -14);
Signal ProductNode_Float2070weight : float ( 5 downto -14 ) := to_float (0.453222,5,14);

Signal ProductNode_Float2070Output_2661: float (5 downto -14);
Signal ProductNode_Float2071weight : float ( 5 downto -14 ) := to_float (0.996146,5,14);

Signal ProductNode_Float2071Output_2662: float (5 downto -14);
Signal SumNode_Float591Output_2663: float (5 downto -14);
Signal ProductNode_Float2072Output_2664: float (5 downto -14);
Signal ProductNode_Float2073weight : float ( 5 downto -14 ) := to_float (0.870697,5,14);

Signal ProductNode_Float2073Output_2665: float (5 downto -14);
Signal ProductNode_Float2074weight : float ( 5 downto -14 ) := to_float (0.753690,5,14);

Signal ProductNode_Float2074Output_2666: float (5 downto -14);
Signal ProductNode_Float2075weight : float ( 5 downto -14 ) := to_float (0.936763,5,14);

Signal ProductNode_Float2075Output_2667: float (5 downto -14);
Signal ProductNode_Float2076weight : float ( 5 downto -14 ) := to_float (0.870404,5,14);

Signal ProductNode_Float2076Output_2668: float (5 downto -14);
Signal ProductNode_Float2077weight : float ( 5 downto -14 ) := to_float (0.933776,5,14);

Signal ProductNode_Float2077Output_2669: float (5 downto -14);
Signal ProductNode_Float2078weight : float ( 5 downto -14 ) := to_float (0.973389,5,14);

Signal ProductNode_Float2078Output_2670: float (5 downto -14);
Signal SumNode_Float592Output_2671: float (5 downto -14);
Signal ProductNode_Float2079Output_2672: float (5 downto -14);
Signal ProductNode_Float2080weight : float ( 5 downto -14 ) := to_float (0.912549,5,14);

Signal ProductNode_Float2080Output_2673: float (5 downto -14);
Signal SumNode_Float593Output_2674: float (5 downto -14);
Signal ProductNode_Float2081Output_2675: float (5 downto -14);
Signal ProductNode_Float2082weight : float ( 5 downto -14 ) := to_float (0.973991,5,14);

Signal ProductNode_Float2082Output_2676: float (5 downto -14);
Signal ProductNode_Float2083weight : float ( 5 downto -14 ) := to_float (0.890735,5,14);

Signal ProductNode_Float2083Output_2677: float (5 downto -14);
Signal ProductNode_Float2084weight : float ( 5 downto -14 ) := to_float (0.382644,5,14);

Signal ProductNode_Float2084Output_2678: float (5 downto -14);
Signal ProductNode_Float2085weight : float ( 5 downto -14 ) := to_float (0.998354,5,14);

Signal ProductNode_Float2085Output_2679: float (5 downto -14);
Signal SumNode_Float594Output_2680: float (5 downto -14);
Signal ProductNode_Float2086Output_2681: float (5 downto -14);
Signal ProductNode_Float2087weight : float ( 5 downto -14 ) := to_float (0.551341,5,14);

Signal ProductNode_Float2087Output_2682: float (5 downto -14);
Signal ProductNode_Float2088weight : float ( 5 downto -14 ) := to_float (0.795357,5,14);

Signal ProductNode_Float2088Output_2683: float (5 downto -14);
Signal ProductNode_Float2089weight : float ( 5 downto -14 ) := to_float (0.948695,5,14);

Signal ProductNode_Float2089Output_2684: float (5 downto -14);
Signal ProductNode_Float2090weight : float ( 5 downto -14 ) := to_float (0.989597,5,14);

Signal ProductNode_Float2090Output_2685: float (5 downto -14);
Signal ProductNode_Float2091weight : float ( 5 downto -14 ) := to_float (0.577708,5,14);

Signal ProductNode_Float2091Output_2686: float (5 downto -14);
Signal ProductNode_Float2092weight : float ( 5 downto -14 ) := to_float (0.981240,5,14);

Signal ProductNode_Float2092Output_2687: float (5 downto -14);
Signal SumNode_Float595Output_2688: float (5 downto -14);
Signal ProductNode_Float2093Output_2689: float (5 downto -14);
Signal ProductNode_Float2094weight : float ( 5 downto -14 ) := to_float (0.712179,5,14);

Signal ProductNode_Float2094Output_2690: float (5 downto -14);
Signal ProductNode_Float2095weight : float ( 5 downto -14 ) := to_float (0.336149,5,14);

Signal ProductNode_Float2095Output_2691: float (5 downto -14);
Signal ProductNode_Float2096weight : float ( 5 downto -14 ) := to_float (0.999140,5,14);

Signal ProductNode_Float2096Output_2692: float (5 downto -14);
Signal SumNode_Float596Output_2693: float (5 downto -14);
Signal ProductNode_Float2097Output_2694: float (5 downto -14);
Signal ProductNode_Float2098weight : float ( 5 downto -14 ) := to_float (0.551341,5,14);

Signal ProductNode_Float2098Output_2695: float (5 downto -14);
Signal ProductNode_Float2099weight : float ( 5 downto -14 ) := to_float (0.926235,5,14);

Signal ProductNode_Float2099Output_2696: float (5 downto -14);
Signal ProductNode_Float2100weight : float ( 5 downto -14 ) := to_float (0.981519,5,14);

Signal ProductNode_Float2100Output_2697: float (5 downto -14);
Signal ProductNode_Float2101weight : float ( 5 downto -14 ) := to_float (0.989597,5,14);

Signal ProductNode_Float2101Output_2698: float (5 downto -14);
Signal ProductNode_Float2102weight : float ( 5 downto -14 ) := to_float (0.986786,5,14);

Signal ProductNode_Float2102Output_2699: float (5 downto -14);
Signal ProductNode_Float2103weight : float ( 5 downto -14 ) := to_float (0.995641,5,14);

Signal ProductNode_Float2103Output_2700: float (5 downto -14);
Signal SumNode_Float597Output_2701: float (5 downto -14);
Signal ProductNode_Float2104Output_2702: float (5 downto -14);
Signal ProductNode_Float2105weight : float ( 5 downto -14 ) := to_float (0.972670,5,14);

Signal ProductNode_Float2105Output_2703: float (5 downto -14);
Signal SumNode_Float598Output_2704: float (5 downto -14);
Signal ProductNode_Float2106Output_2705: float (5 downto -14);
Signal ProductNode_Float2107weight : float ( 5 downto -14 ) := to_float (0.991382,5,14);

Signal ProductNode_Float2107Output_2706: float (5 downto -14);
Signal SumNode_Float599Output_2707: float (5 downto -14);
Signal ProductNode_Float2108Output_2708: float (5 downto -14);
Signal ProductNode_Float2109weight : float ( 5 downto -14 ) := to_float (0.987767,5,14);

Signal ProductNode_Float2109Output_2709: float (5 downto -14);
Signal SumNode_Float600Output_2710: float (5 downto -14);
Signal ProductNode_Float2110Output_2711: float (5 downto -14);
Signal ProductNode_Float2111weight : float ( 5 downto -14 ) := to_float (0.965849,5,14);

Signal ProductNode_Float2111Output_2712: float (5 downto -14);
Signal ProductNode_Float2112weight : float ( 5 downto -14 ) := to_float (0.692695,5,14);

Signal ProductNode_Float2112Output_2713: float (5 downto -14);
Signal SumNode_Float601Output_2714: float (5 downto -14);
Signal ProductNode_Float2113Output_2715: float (5 downto -14);
Signal ProductNode_Float2114weight : float ( 5 downto -14 ) := to_float (0.880399,5,14);

Signal ProductNode_Float2114Output_2716: float (5 downto -14);
Signal ProductNode_Float2115weight : float ( 5 downto -14 ) := to_float (0.997554,5,14);

Signal ProductNode_Float2115Output_2717: float (5 downto -14);
Signal ProductNode_Float2116weight : float ( 5 downto -14 ) := to_float (0.414069,5,14);

Signal ProductNode_Float2116Output_2718: float (5 downto -14);
Signal SumNode_Float602Output_2719: float (5 downto -14);
Signal ProductNode_Float2117Output_2720: float (5 downto -14);
Signal ProductNode_Float2118weight : float ( 5 downto -14 ) := to_float (0.919660,5,14);

Signal ProductNode_Float2118Output_2721: float (5 downto -14);
Signal ProductNode_Float2119weight : float ( 5 downto -14 ) := to_float (0.806938,5,14);

Signal ProductNode_Float2119Output_2722: float (5 downto -14);
Signal SumNode_Float603Output_2723: float (5 downto -14);
Signal ProductNode_Float2120Output_2724: float (5 downto -14);
Signal ProductNode_Float2121weight : float ( 5 downto -14 ) := to_float (0.860235,5,14);

Signal ProductNode_Float2121Output_2725: float (5 downto -14);
Signal ProductNode_Float2122weight : float ( 5 downto -14 ) := to_float (0.989739,5,14);

Signal ProductNode_Float2122Output_2726: float (5 downto -14);
Signal ProductNode_Float2123weight : float ( 5 downto -14 ) := to_float (0.549861,5,14);

Signal ProductNode_Float2123Output_2727: float (5 downto -14);
Signal SumNode_Float604Output_2728: float (5 downto -14);
Signal ProductNode_Float2124Output_2729: float (5 downto -14);
Signal SumNode_Float605Output_2730: float (5 downto -14);
Signal ProductNode_Float2125Output_2731: float (5 downto -14);
Signal ProductNode_Float2126weight : float ( 5 downto -14 ) := to_float (0.984104,5,14);

Signal ProductNode_Float2126Output_2732: float (5 downto -14);
Signal ProductNode_Float2127weight : float ( 5 downto -14 ) := to_float (0.793165,5,14);

Signal ProductNode_Float2127Output_2733: float (5 downto -14);
Signal ProductNode_Float2128weight : float ( 5 downto -14 ) := to_float (0.927417,5,14);

Signal ProductNode_Float2128Output_2734: float (5 downto -14);
Signal SumNode_Float606Output_2735: float (5 downto -14);
Signal ProductNode_Float2129Output_2736: float (5 downto -14);
Signal ProductNode_Float2130weight : float ( 5 downto -14 ) := to_float (0.726095,5,14);

Signal ProductNode_Float2130Output_2737: float (5 downto -14);
Signal ProductNode_Float2131weight : float ( 5 downto -14 ) := to_float (0.988880,5,14);

Signal ProductNode_Float2131Output_2738: float (5 downto -14);
Signal ProductNode_Float2132weight : float ( 5 downto -14 ) := to_float (0.558577,5,14);

Signal ProductNode_Float2132Output_2739: float (5 downto -14);
Signal SumNode_Float607Output_2740: float (5 downto -14);
Signal ProductNode_Float2133Output_2741: float (5 downto -14);
Signal ProductNode_Float2134weight : float ( 5 downto -14 ) := to_float (0.649155,5,14);

Signal ProductNode_Float2134Output_2742: float (5 downto -14);
Signal ProductNode_Float2135weight : float ( 5 downto -14 ) := to_float (0.975801,5,14);

Signal ProductNode_Float2135Output_2743: float (5 downto -14);
Signal SumNode_Float608Output_2744: float (5 downto -14);
Signal ProductNode_Float2136Output_2745: float (5 downto -14);
Signal ProductNode_Float2137weight : float ( 5 downto -14 ) := to_float (0.955917,5,14);

Signal ProductNode_Float2137Output_2746: float (5 downto -14);
Signal ProductNode_Float2138weight : float ( 5 downto -14 ) := to_float (0.985013,5,14);

Signal ProductNode_Float2138Output_2747: float (5 downto -14);
Signal ProductNode_Float2139weight : float ( 5 downto -14 ) := to_float (0.592017,5,14);

Signal ProductNode_Float2139Output_2748: float (5 downto -14);
Signal SumNode_Float609Output_2749: float (5 downto -14);
Signal ProductNode_Float2140Output_2750: float (5 downto -14);
Signal SumNode_Float610Output_2751: float (5 downto -14);
Signal ProductNode_Float2141Output_2752: float (5 downto -14);
Signal ProductNode_Float2142weight : float ( 5 downto -14 ) := to_float (0.598812,5,14);

Signal ProductNode_Float2142Output_2753: float (5 downto -14);
Signal SumNode_Float611Output_2754: float (5 downto -14);
Signal ProductNode_Float2143Output_2755: float (5 downto -14);
Signal ProductNode_Float2144weight : float ( 5 downto -14 ) := to_float (0.807423,5,14);

Signal ProductNode_Float2144Output_2756: float (5 downto -14);
Signal ProductNode_Float2145weight : float ( 5 downto -14 ) := to_float (0.919372,5,14);

Signal ProductNode_Float2145Output_2757: float (5 downto -14);
Signal SumNode_Float612Output_2758: float (5 downto -14);
Signal ProductNode_Float2146Output_2759: float (5 downto -14);
Signal ProductNode_Float2147weight : float ( 5 downto -14 ) := to_float (0.694473,5,14);

Signal ProductNode_Float2147Output_2760: float (5 downto -14);
Signal ProductNode_Float2148weight : float ( 5 downto -14 ) := to_float (0.843444,5,14);

Signal ProductNode_Float2148Output_2761: float (5 downto -14);
Signal ProductNode_Float2149weight : float ( 5 downto -14 ) := to_float (0.682797,5,14);

Signal ProductNode_Float2149Output_2762: float (5 downto -14);
Signal ProductNode_Float2150weight : float ( 5 downto -14 ) := to_float (0.968381,5,14);

Signal ProductNode_Float2150Output_2763: float (5 downto -14);
Signal SumNode_Float613Output_2764: float (5 downto -14);
Signal ProductNode_Float2151Output_2765: float (5 downto -14);
Signal ProductNode_Float2152weight : float ( 5 downto -14 ) := to_float (0.965376,5,14);

Signal ProductNode_Float2152Output_2766: float (5 downto -14);
Signal ProductNode_Float2153weight : float ( 5 downto -14 ) := to_float (0.697447,5,14);

Signal ProductNode_Float2153Output_2767: float (5 downto -14);
Signal SumNode_Float614Output_2768: float (5 downto -14);
Signal ProductNode_Float2154Output_2769: float (5 downto -14);
Signal ProductNode_Float2155weight : float ( 5 downto -14 ) := to_float (0.965849,5,14);

Signal ProductNode_Float2155Output_2770: float (5 downto -14);
Signal ProductNode_Float2156weight : float ( 5 downto -14 ) := to_float (0.692695,5,14);

Signal ProductNode_Float2156Output_2771: float (5 downto -14);
Signal SumNode_Float615Output_2772: float (5 downto -14);
Signal ProductNode_Float2157Output_2773: float (5 downto -14);
Signal ProductNode_Float2158weight : float ( 5 downto -14 ) := to_float (0.880399,5,14);

Signal ProductNode_Float2158Output_2774: float (5 downto -14);
Signal ProductNode_Float2159weight : float ( 5 downto -14 ) := to_float (0.997554,5,14);

Signal ProductNode_Float2159Output_2775: float (5 downto -14);
Signal ProductNode_Float2160weight : float ( 5 downto -14 ) := to_float (0.414069,5,14);

Signal ProductNode_Float2160Output_2776: float (5 downto -14);
Signal SumNode_Float616Output_2777: float (5 downto -14);
Signal ProductNode_Float2161Output_2778: float (5 downto -14);
Signal ProductNode_Float2162weight : float ( 5 downto -14 ) := to_float (0.919660,5,14);

Signal ProductNode_Float2162Output_2779: float (5 downto -14);
Signal ProductNode_Float2163weight : float ( 5 downto -14 ) := to_float (0.806938,5,14);

Signal ProductNode_Float2163Output_2780: float (5 downto -14);
Signal SumNode_Float617Output_2781: float (5 downto -14);
Signal ProductNode_Float2164Output_2782: float (5 downto -14);
Signal ProductNode_Float2165weight : float ( 5 downto -14 ) := to_float (0.860235,5,14);

Signal ProductNode_Float2165Output_2783: float (5 downto -14);
Signal ProductNode_Float2166weight : float ( 5 downto -14 ) := to_float (0.989739,5,14);

Signal ProductNode_Float2166Output_2784: float (5 downto -14);
Signal ProductNode_Float2167weight : float ( 5 downto -14 ) := to_float (0.549861,5,14);

Signal ProductNode_Float2167Output_2785: float (5 downto -14);
Signal SumNode_Float618Output_2786: float (5 downto -14);
Signal ProductNode_Float2168Output_2787: float (5 downto -14);
Signal SumNode_Float619Output_2788: float (5 downto -14);
Signal ProductNode_Float2169Output_2789: float (5 downto -14);
Signal ProductNode_Float2170weight : float ( 5 downto -14 ) := to_float (0.932937,5,14);

Signal ProductNode_Float2170Output_2790: float (5 downto -14);
Signal ProductNode_Float2171weight : float ( 5 downto -14 ) := to_float (0.793165,5,14);

Signal ProductNode_Float2171Output_2791: float (5 downto -14);
Signal ProductNode_Float2172weight : float ( 5 downto -14 ) := to_float (0.927417,5,14);

Signal ProductNode_Float2172Output_2792: float (5 downto -14);
Signal SumNode_Float620Output_2793: float (5 downto -14);
Signal ProductNode_Float2173Output_2794: float (5 downto -14);
Signal ProductNode_Float2174weight : float ( 5 downto -14 ) := to_float (0.726095,5,14);

Signal ProductNode_Float2174Output_2795: float (5 downto -14);
Signal ProductNode_Float2175weight : float ( 5 downto -14 ) := to_float (0.988880,5,14);

Signal ProductNode_Float2175Output_2796: float (5 downto -14);
Signal ProductNode_Float2176weight : float ( 5 downto -14 ) := to_float (0.558577,5,14);

Signal ProductNode_Float2176Output_2797: float (5 downto -14);
Signal SumNode_Float621Output_2798: float (5 downto -14);
Signal ProductNode_Float2177Output_2799: float (5 downto -14);
Signal ProductNode_Float2178weight : float ( 5 downto -14 ) := to_float (0.649155,5,14);

Signal ProductNode_Float2178Output_2800: float (5 downto -14);
Signal ProductNode_Float2179weight : float ( 5 downto -14 ) := to_float (0.975801,5,14);

Signal ProductNode_Float2179Output_2801: float (5 downto -14);
Signal SumNode_Float622Output_2802: float (5 downto -14);
Signal ProductNode_Float2180Output_2803: float (5 downto -14);
Signal ProductNode_Float2181weight : float ( 5 downto -14 ) := to_float (0.955917,5,14);

Signal ProductNode_Float2181Output_2804: float (5 downto -14);
Signal ProductNode_Float2182weight : float ( 5 downto -14 ) := to_float (0.985013,5,14);

Signal ProductNode_Float2182Output_2805: float (5 downto -14);
Signal ProductNode_Float2183weight : float ( 5 downto -14 ) := to_float (0.592017,5,14);

Signal ProductNode_Float2183Output_2806: float (5 downto -14);
Signal SumNode_Float623Output_2807: float (5 downto -14);
Signal ProductNode_Float2184Output_2808: float (5 downto -14);
Signal SumNode_Float624Output_2809: float (5 downto -14);
Signal ProductNode_Float2185Output_2810: float (5 downto -14);
Signal ProductNode_Float2186weight : float ( 5 downto -14 ) := to_float (0.782438,5,14);

Signal ProductNode_Float2186Output_2811: float (5 downto -14);
Signal SumNode_Float625Output_2812: float (5 downto -14);
Signal ProductNode_Float2187Output_2813: float (5 downto -14);
Signal ProductNode_Float2188weight : float ( 5 downto -14 ) := to_float (0.623360,5,14);

Signal ProductNode_Float2188Output_2814: float (5 downto -14);
Signal ProductNode_Float2189weight : float ( 5 downto -14 ) := to_float (0.980424,5,14);

Signal ProductNode_Float2189Output_2815: float (5 downto -14);
Signal SumNode_Float626Output_2816: float (5 downto -14);
Signal ProductNode_Float2190Output_2817: float (5 downto -14);
Signal ProductNode_Float2191weight : float ( 5 downto -14 ) := to_float (0.694473,5,14);

Signal ProductNode_Float2191Output_2818: float (5 downto -14);
Signal ProductNode_Float2192weight : float ( 5 downto -14 ) := to_float (0.894649,5,14);

Signal ProductNode_Float2192Output_2819: float (5 downto -14);
Signal ProductNode_Float2193weight : float ( 5 downto -14 ) := to_float (0.482891,5,14);

Signal ProductNode_Float2193Output_2820: float (5 downto -14);
Signal ProductNode_Float2194weight : float ( 5 downto -14 ) := to_float (0.994693,5,14);

Signal ProductNode_Float2194Output_2821: float (5 downto -14);
Signal SumNode_Float627Output_2822: float (5 downto -14);
Signal ProductNode_Float2195Output_2823: float (5 downto -14);
Signal ProductNode_Float2196weight : float ( 5 downto -14 ) := to_float (0.965376,5,14);

Signal ProductNode_Float2196Output_2824: float (5 downto -14);
Signal ProductNode_Float2197weight : float ( 5 downto -14 ) := to_float (0.964572,5,14);

Signal ProductNode_Float2197Output_2825: float (5 downto -14);
Signal SumNode_Float628Output_2826: float (5 downto -14);
Signal ProductNode_Float2198Output_2827: float (5 downto -14);
Signal SumNode_Float629Output_2828: float (5 downto -14);
Signal ProductNode_Float2199Output_2829: float (5 downto -14);
Signal ProductNode_Float2200weight : float ( 5 downto -14 ) := to_float (0.625034,5,14);

Signal ProductNode_Float2200Output_2830: float (5 downto -14);
Signal ProductNode_Float2201weight : float ( 5 downto -14 ) := to_float (0.965849,5,14);

Signal ProductNode_Float2201Output_2831: float (5 downto -14);
Signal ProductNode_Float2202weight : float ( 5 downto -14 ) := to_float (0.692695,5,14);

Signal ProductNode_Float2202Output_2832: float (5 downto -14);
Signal SumNode_Float630Output_2833: float (5 downto -14);
Signal ProductNode_Float2203Output_2834: float (5 downto -14);
Signal ProductNode_Float2204weight : float ( 5 downto -14 ) := to_float (0.880399,5,14);

Signal ProductNode_Float2204Output_2835: float (5 downto -14);
Signal ProductNode_Float2205weight : float ( 5 downto -14 ) := to_float (0.966381,5,14);

Signal ProductNode_Float2205Output_2836: float (5 downto -14);
Signal ProductNode_Float2206weight : float ( 5 downto -14 ) := to_float (0.690672,5,14);

Signal ProductNode_Float2206Output_2837: float (5 downto -14);
Signal SumNode_Float631Output_2838: float (5 downto -14);
Signal ProductNode_Float2207Output_2839: float (5 downto -14);
Signal ProductNode_Float2208weight : float ( 5 downto -14 ) := to_float (0.919660,5,14);

Signal ProductNode_Float2208Output_2840: float (5 downto -14);
Signal ProductNode_Float2209weight : float ( 5 downto -14 ) := to_float (0.806938,5,14);

Signal ProductNode_Float2209Output_2841: float (5 downto -14);
Signal SumNode_Float632Output_2842: float (5 downto -14);
Signal ProductNode_Float2210Output_2843: float (5 downto -14);
Signal ProductNode_Float2211weight : float ( 5 downto -14 ) := to_float (0.860235,5,14);

Signal ProductNode_Float2211Output_2844: float (5 downto -14);
Signal ProductNode_Float2212weight : float ( 5 downto -14 ) := to_float (0.941870,5,14);

Signal ProductNode_Float2212Output_2845: float (5 downto -14);
Signal ProductNode_Float2213weight : float ( 5 downto -14 ) := to_float (0.763101,5,14);

Signal ProductNode_Float2213Output_2846: float (5 downto -14);
Signal SumNode_Float633Output_2847: float (5 downto -14);
Signal ProductNode_Float2214Output_2848: float (5 downto -14);
Signal SumNode_Float634Output_2849: float (5 downto -14);
Signal ProductNode_Float2215Output_2850: float (5 downto -14);
Signal ProductNode_Float2216weight : float ( 5 downto -14 ) := to_float (0.924413,5,14);

Signal ProductNode_Float2216Output_2851: float (5 downto -14);
Signal ProductNode_Float2217weight : float ( 5 downto -14 ) := to_float (0.793165,5,14);

Signal ProductNode_Float2217Output_2852: float (5 downto -14);
Signal ProductNode_Float2218weight : float ( 5 downto -14 ) := to_float (0.927417,5,14);

Signal ProductNode_Float2218Output_2853: float (5 downto -14);
Signal SumNode_Float635Output_2854: float (5 downto -14);
Signal ProductNode_Float2219Output_2855: float (5 downto -14);
Signal ProductNode_Float2220weight : float ( 5 downto -14 ) := to_float (0.726095,5,14);

Signal ProductNode_Float2220Output_2856: float (5 downto -14);
Signal ProductNode_Float2221weight : float ( 5 downto -14 ) := to_float (0.909585,5,14);

Signal ProductNode_Float2221Output_2857: float (5 downto -14);
Signal ProductNode_Float2222weight : float ( 5 downto -14 ) := to_float (0.822920,5,14);

Signal ProductNode_Float2222Output_2858: float (5 downto -14);
Signal SumNode_Float636Output_2859: float (5 downto -14);
Signal ProductNode_Float2223Output_2860: float (5 downto -14);
Signal ProductNode_Float2224weight : float ( 5 downto -14 ) := to_float (0.649155,5,14);

Signal ProductNode_Float2224Output_2861: float (5 downto -14);
Signal ProductNode_Float2225weight : float ( 5 downto -14 ) := to_float (0.975801,5,14);

Signal ProductNode_Float2225Output_2862: float (5 downto -14);
Signal SumNode_Float637Output_2863: float (5 downto -14);
Signal ProductNode_Float2226Output_2864: float (5 downto -14);
Signal ProductNode_Float2227weight : float ( 5 downto -14 ) := to_float (0.955917,5,14);

Signal ProductNode_Float2227Output_2865: float (5 downto -14);
Signal ProductNode_Float2228weight : float ( 5 downto -14 ) := to_float (0.790147,5,14);

Signal ProductNode_Float2228Output_2866: float (5 downto -14);
Signal ProductNode_Float2229weight : float ( 5 downto -14 ) := to_float (0.929014,5,14);

Signal ProductNode_Float2229Output_2867: float (5 downto -14);
Signal SumNode_Float638Output_2868: float (5 downto -14);
Signal ProductNode_Float2230Output_2869: float (5 downto -14);
Signal SumNode_Float639Output_2870: float (5 downto -14);
Signal ProductNode_Float2231Output_2871: float (5 downto -14);
Signal ProductNode_Float2232weight : float ( 5 downto -14 ) := to_float (0.798666,5,14);

Signal ProductNode_Float2232Output_2872: float (5 downto -14);
Signal SumNode_Float640Output_2873: float (5 downto -14);
Signal ProductNode_Float2233Output_2874: float (5 downto -14);
Signal ProductNode_Float2234weight : float ( 5 downto -14 ) := to_float (0.807423,5,14);

Signal ProductNode_Float2234Output_2875: float (5 downto -14);
Signal ProductNode_Float2235weight : float ( 5 downto -14 ) := to_float (0.919372,5,14);

Signal ProductNode_Float2235Output_2876: float (5 downto -14);
Signal SumNode_Float641Output_2877: float (5 downto -14);
Signal ProductNode_Float2236Output_2878: float (5 downto -14);
Signal ProductNode_Float2237weight : float ( 5 downto -14 ) := to_float (0.579487,5,14);

Signal ProductNode_Float2237Output_2879: float (5 downto -14);
Signal ProductNode_Float2238weight : float ( 5 downto -14 ) := to_float (0.790558,5,14);

Signal ProductNode_Float2238Output_2880: float (5 downto -14);
Signal ProductNode_Float2239weight : float ( 5 downto -14 ) := to_float (0.682797,5,14);

Signal ProductNode_Float2239Output_2881: float (5 downto -14);
Signal ProductNode_Float2240weight : float ( 5 downto -14 ) := to_float (0.968381,5,14);

Signal ProductNode_Float2240Output_2882: float (5 downto -14);
Signal SumNode_Float642Output_2883: float (5 downto -14);
Signal ProductNode_Float2241Output_2884: float (5 downto -14);
Signal ProductNode_Float2242weight : float ( 5 downto -14 ) := to_float (0.986575,5,14);

Signal ProductNode_Float2242Output_2885: float (5 downto -14);
Signal ProductNode_Float2243weight : float ( 5 downto -14 ) := to_float (0.578242,5,14);

Signal ProductNode_Float2243Output_2886: float (5 downto -14);
Signal SumNode_Float643Output_2887: float (5 downto -14);
Signal ProductNode_Float2244Output_2888: float (5 downto -14);
Signal ProductNode_Float2245weight : float ( 5 downto -14 ) := to_float (0.965849,5,14);

Signal ProductNode_Float2245Output_2889: float (5 downto -14);
Signal ProductNode_Float2246weight : float ( 5 downto -14 ) := to_float (0.692695,5,14);

Signal ProductNode_Float2246Output_2890: float (5 downto -14);
Signal SumNode_Float644Output_2891: float (5 downto -14);
Signal ProductNode_Float2247Output_2892: float (5 downto -14);
Signal ProductNode_Float2248weight : float ( 5 downto -14 ) := to_float (0.880399,5,14);

Signal ProductNode_Float2248Output_2893: float (5 downto -14);
Signal ProductNode_Float2249weight : float ( 5 downto -14 ) := to_float (0.966381,5,14);

Signal ProductNode_Float2249Output_2894: float (5 downto -14);
Signal ProductNode_Float2250weight : float ( 5 downto -14 ) := to_float (0.690672,5,14);

Signal ProductNode_Float2250Output_2895: float (5 downto -14);
Signal SumNode_Float645Output_2896: float (5 downto -14);
Signal ProductNode_Float2251Output_2897: float (5 downto -14);
Signal ProductNode_Float2252weight : float ( 5 downto -14 ) := to_float (0.919660,5,14);

Signal ProductNode_Float2252Output_2898: float (5 downto -14);
Signal ProductNode_Float2253weight : float ( 5 downto -14 ) := to_float (0.806938,5,14);

Signal ProductNode_Float2253Output_2899: float (5 downto -14);
Signal SumNode_Float646Output_2900: float (5 downto -14);
Signal ProductNode_Float2254Output_2901: float (5 downto -14);
Signal ProductNode_Float2255weight : float ( 5 downto -14 ) := to_float (0.860235,5,14);

Signal ProductNode_Float2255Output_2902: float (5 downto -14);
Signal ProductNode_Float2256weight : float ( 5 downto -14 ) := to_float (0.941870,5,14);

Signal ProductNode_Float2256Output_2903: float (5 downto -14);
Signal ProductNode_Float2257weight : float ( 5 downto -14 ) := to_float (0.763101,5,14);

Signal ProductNode_Float2257Output_2904: float (5 downto -14);
Signal SumNode_Float647Output_2905: float (5 downto -14);
Signal ProductNode_Float2258Output_2906: float (5 downto -14);
Signal SumNode_Float648Output_2907: float (5 downto -14);
Signal ProductNode_Float2259Output_2908: float (5 downto -14);
Signal ProductNode_Float2260weight : float ( 5 downto -14 ) := to_float (0.693688,5,14);

Signal ProductNode_Float2260Output_2909: float (5 downto -14);
Signal ProductNode_Float2261weight : float ( 5 downto -14 ) := to_float (0.793165,5,14);

Signal ProductNode_Float2261Output_2910: float (5 downto -14);
Signal ProductNode_Float2262weight : float ( 5 downto -14 ) := to_float (0.927417,5,14);

Signal ProductNode_Float2262Output_2911: float (5 downto -14);
Signal SumNode_Float649Output_2912: float (5 downto -14);
Signal ProductNode_Float2263Output_2913: float (5 downto -14);
Signal ProductNode_Float2264weight : float ( 5 downto -14 ) := to_float (0.726095,5,14);

Signal ProductNode_Float2264Output_2914: float (5 downto -14);
Signal ProductNode_Float2265weight : float ( 5 downto -14 ) := to_float (0.909585,5,14);

Signal ProductNode_Float2265Output_2915: float (5 downto -14);
Signal ProductNode_Float2266weight : float ( 5 downto -14 ) := to_float (0.822920,5,14);

Signal ProductNode_Float2266Output_2916: float (5 downto -14);
Signal SumNode_Float650Output_2917: float (5 downto -14);
Signal ProductNode_Float2267Output_2918: float (5 downto -14);
Signal ProductNode_Float2268weight : float ( 5 downto -14 ) := to_float (0.649155,5,14);

Signal ProductNode_Float2268Output_2919: float (5 downto -14);
Signal ProductNode_Float2269weight : float ( 5 downto -14 ) := to_float (0.975801,5,14);

Signal ProductNode_Float2269Output_2920: float (5 downto -14);
Signal SumNode_Float651Output_2921: float (5 downto -14);
Signal ProductNode_Float2270Output_2922: float (5 downto -14);
Signal ProductNode_Float2271weight : float ( 5 downto -14 ) := to_float (0.955917,5,14);

Signal ProductNode_Float2271Output_2923: float (5 downto -14);
Signal ProductNode_Float2272weight : float ( 5 downto -14 ) := to_float (0.790147,5,14);

Signal ProductNode_Float2272Output_2924: float (5 downto -14);
Signal ProductNode_Float2273weight : float ( 5 downto -14 ) := to_float (0.929014,5,14);

Signal ProductNode_Float2273Output_2925: float (5 downto -14);
Signal SumNode_Float652Output_2926: float (5 downto -14);
Signal ProductNode_Float2274Output_2927: float (5 downto -14);
Signal SumNode_Float653Output_2928: float (5 downto -14);
Signal ProductNode_Float2275Output_2929: float (5 downto -14);
Signal ProductNode_Float2276weight : float ( 5 downto -14 ) := to_float (0.965586,5,14);

Signal ProductNode_Float2276Output_2930: float (5 downto -14);
Signal SumNode_Float654Output_2931: float (5 downto -14);
Signal ProductNode_Float2277Output_2932: float (5 downto -14);
Signal ProductNode_Float2278weight : float ( 5 downto -14 ) := to_float (0.623360,5,14);

Signal ProductNode_Float2278Output_2933: float (5 downto -14);
Signal ProductNode_Float2279weight : float ( 5 downto -14 ) := to_float (0.980424,5,14);

Signal ProductNode_Float2279Output_2934: float (5 downto -14);
Signal SumNode_Float655Output_2935: float (5 downto -14);
Signal ProductNode_Float2280Output_2936: float (5 downto -14);
Signal ProductNode_Float2281weight : float ( 5 downto -14 ) := to_float (0.579487,5,14);

Signal ProductNode_Float2281Output_2937: float (5 downto -14);
Signal ProductNode_Float2282weight : float ( 5 downto -14 ) := to_float (0.928799,5,14);

Signal ProductNode_Float2282Output_2938: float (5 downto -14);
Signal ProductNode_Float2283weight : float ( 5 downto -14 ) := to_float (0.482891,5,14);

Signal ProductNode_Float2283Output_2939: float (5 downto -14);
Signal ProductNode_Float2284weight : float ( 5 downto -14 ) := to_float (0.994693,5,14);

Signal ProductNode_Float2284Output_2940: float (5 downto -14);
Signal SumNode_Float656Output_2941: float (5 downto -14);
Signal ProductNode_Float2285Output_2942: float (5 downto -14);
Signal ProductNode_Float2286weight : float ( 5 downto -14 ) := to_float (0.986575,5,14);

Signal ProductNode_Float2286Output_2943: float (5 downto -14);
Signal ProductNode_Float2287weight : float ( 5 downto -14 ) := to_float (0.986723,5,14);

Signal ProductNode_Float2287Output_2944: float (5 downto -14);
Signal SumNode_Float657Output_2945: float (5 downto -14);
Signal ProductNode_Float2288Output_2946: float (5 downto -14);
Signal SumNode_Float658Output_2947: float (5 downto -14);
Signal ProductNode_Float2289Output_2948: float (5 downto -14);
Signal ProductNode_Float2290weight : float ( 5 downto -14 ) := to_float (0.980149,5,14);

Signal ProductNode_Float2290Output_2949: float (5 downto -14);
Signal SumNode_Float659Output_2950: float (5 downto -14);
Signal ProductNode_Float2291Output_2951: float (5 downto -14);
Signal SumNode_Float660Output_2952: float (5 downto -14);
Signal ProductNode_Float2292Output_2953: float (5 downto -14);
Signal SumNode_Float661Output_2954: float (5 downto -14);
Signal ProductNode_Float2293Output_2955: float (5 downto -14);
Signal SumNode_Float662Output_2956: float (5 downto -14);

 
begin 
ProductNode_Float0: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float0weight,v4,ProductNode_Float0Output_0);

ProductNode_Float1: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1weight,v8,ProductNode_Float1Output_1);

ProductNode_Float2: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2weight,vb8,ProductNode_Float2Output_2);

SumNode_Float0: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2Output_2,ProductNode_Float1Output_1,SumNode_Float0Output_3);

ProductNode_Float3: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v7,SumNode_Float0Output_3,ProductNode_Float3Output_4);

ProductNode_Float4: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float4weight,v3,ProductNode_Float4Output_5);

ProductNode_Float5: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float5weight,ProductNode_Float4Output_5,ProductNode_Float5Output_6);

ProductNode_Float6: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float6weight,ProductNode_Float5Output_6,ProductNode_Float6Output_7);

ProductNode_Float7: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float7weight,vb3,ProductNode_Float7Output_8);

ProductNode_Float8: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float8weight,ProductNode_Float7Output_8,ProductNode_Float8Output_9);

ProductNode_Float9: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float9weight,ProductNode_Float8Output_9,ProductNode_Float9Output_10);

SumNode_Float1: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float9Output_10,ProductNode_Float6Output_7,SumNode_Float1Output_11);

ProductNode_Float10: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float1Output_11,ProductNode_Float3Output_4,ProductNode_Float10Output_12);

ProductNode_Float11: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float11weight,ProductNode_Float10Output_12,ProductNode_Float11Output_13);

ProductNode_Float12: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float12weight,v8,ProductNode_Float12Output_14);

ProductNode_Float13: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float13weight,vb8,ProductNode_Float13Output_15);

SumNode_Float2: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float13Output_15,ProductNode_Float12Output_14,SumNode_Float2Output_16);

ProductNode_Float14: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb7,SumNode_Float2Output_16,ProductNode_Float14Output_17);

ProductNode_Float15: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float15weight,v3,ProductNode_Float15Output_18);

ProductNode_Float16: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float16weight,ProductNode_Float4Output_5,ProductNode_Float16Output_19);

ProductNode_Float17: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float17weight,ProductNode_Float16Output_19,ProductNode_Float17Output_20);

ProductNode_Float18: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float18weight,vb3,ProductNode_Float18Output_21);

ProductNode_Float19: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float19weight,ProductNode_Float7Output_8,ProductNode_Float19Output_22);

ProductNode_Float20: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float20weight,ProductNode_Float19Output_22,ProductNode_Float20Output_23);

SumNode_Float3: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float20Output_23,ProductNode_Float17Output_20,SumNode_Float3Output_24);

ProductNode_Float21: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float3Output_24,ProductNode_Float14Output_17,ProductNode_Float21Output_25);

ProductNode_Float22: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float22weight,ProductNode_Float21Output_25,ProductNode_Float22Output_26);

SumNode_Float4: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float22Output_26,ProductNode_Float11Output_13,SumNode_Float4Output_27);

ProductNode_Float23: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float4Output_27,ProductNode_Float0Output_0,ProductNode_Float23Output_28);

ProductNode_Float24: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float24weight,ProductNode_Float23Output_28,ProductNode_Float24Output_29);

ProductNode_Float25: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float25weight,vb4,ProductNode_Float25Output_30);

ProductNode_Float26: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float26weight,v8,ProductNode_Float26Output_31);

ProductNode_Float27: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float27weight,vb8,ProductNode_Float27Output_32);

SumNode_Float5: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float27Output_32,ProductNode_Float26Output_31,SumNode_Float5Output_33);

ProductNode_Float28: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v7,SumNode_Float5Output_33,ProductNode_Float28Output_34);

ProductNode_Float29: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float29weight,v3,ProductNode_Float29Output_35);

ProductNode_Float30: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float30weight,ProductNode_Float29Output_35,ProductNode_Float30Output_36);

ProductNode_Float31: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float31weight,ProductNode_Float30Output_36,ProductNode_Float31Output_37);

ProductNode_Float32: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float32weight,vb3,ProductNode_Float32Output_38);

ProductNode_Float33: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float33weight,ProductNode_Float32Output_38,ProductNode_Float33Output_39);

ProductNode_Float34: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float34weight,ProductNode_Float33Output_39,ProductNode_Float34Output_40);

SumNode_Float6: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float34Output_40,ProductNode_Float31Output_37,SumNode_Float6Output_41);

ProductNode_Float35: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float6Output_41,ProductNode_Float28Output_34,ProductNode_Float35Output_42);

ProductNode_Float36: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float36weight,ProductNode_Float35Output_42,ProductNode_Float36Output_43);

ProductNode_Float37: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float37weight,v8,ProductNode_Float37Output_44);

ProductNode_Float38: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float38weight,vb8,ProductNode_Float38Output_45);

SumNode_Float7: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float38Output_45,ProductNode_Float37Output_44,SumNode_Float7Output_46);

ProductNode_Float39: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb7,SumNode_Float7Output_46,ProductNode_Float39Output_47);

ProductNode_Float40: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float40weight,v3,ProductNode_Float40Output_48);

ProductNode_Float41: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float41weight,ProductNode_Float29Output_35,ProductNode_Float41Output_49);

ProductNode_Float42: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float42weight,ProductNode_Float41Output_49,ProductNode_Float42Output_50);

ProductNode_Float43: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float43weight,vb3,ProductNode_Float43Output_51);

ProductNode_Float44: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float44weight,ProductNode_Float32Output_38,ProductNode_Float44Output_52);

ProductNode_Float45: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float45weight,ProductNode_Float44Output_52,ProductNode_Float45Output_53);

SumNode_Float8: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float45Output_53,ProductNode_Float42Output_50,SumNode_Float8Output_54);

ProductNode_Float46: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float8Output_54,ProductNode_Float39Output_47,ProductNode_Float46Output_55);

ProductNode_Float47: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float47weight,ProductNode_Float46Output_55,ProductNode_Float47Output_56);

SumNode_Float9: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float47Output_56,ProductNode_Float36Output_43,SumNode_Float9Output_57);

ProductNode_Float48: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float9Output_57,ProductNode_Float25Output_30,ProductNode_Float48Output_58);

ProductNode_Float49: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float49weight,ProductNode_Float48Output_58,ProductNode_Float49Output_59);

SumNode_Float10: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float49Output_59,ProductNode_Float24Output_29,SumNode_Float10Output_60);

ProductNode_Float50: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v5,SumNode_Float10Output_60,ProductNode_Float50Output_61);

ProductNode_Float51: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float51weight,ProductNode_Float50Output_61,ProductNode_Float51Output_62);

ProductNode_Float52: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float52weight,v4,ProductNode_Float52Output_63);

ProductNode_Float53: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float53weight,v8,ProductNode_Float53Output_64);

ProductNode_Float54: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float54weight,vb8,ProductNode_Float54Output_65);

SumNode_Float11: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float54Output_65,ProductNode_Float53Output_64,SumNode_Float11Output_66);

ProductNode_Float55: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v7,SumNode_Float11Output_66,ProductNode_Float55Output_67);

ProductNode_Float56: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float56weight,v3,ProductNode_Float56Output_68);

ProductNode_Float57: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float57weight,ProductNode_Float4Output_5,ProductNode_Float57Output_69);

ProductNode_Float58: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float58weight,ProductNode_Float5Output_6,ProductNode_Float58Output_70);

ProductNode_Float59: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float59weight,vb3,ProductNode_Float59Output_71);

ProductNode_Float60: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float60weight,ProductNode_Float7Output_8,ProductNode_Float60Output_72);

ProductNode_Float61: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float61weight,ProductNode_Float8Output_9,ProductNode_Float61Output_73);

SumNode_Float12: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float61Output_73,ProductNode_Float58Output_70,SumNode_Float12Output_74);

ProductNode_Float62: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float12Output_74,ProductNode_Float55Output_67,ProductNode_Float62Output_75);

ProductNode_Float63: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float63weight,ProductNode_Float62Output_75,ProductNode_Float63Output_76);

ProductNode_Float64: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float64weight,v8,ProductNode_Float64Output_77);

ProductNode_Float65: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float65weight,vb8,ProductNode_Float65Output_78);

SumNode_Float13: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float65Output_78,ProductNode_Float64Output_77,SumNode_Float13Output_79);

ProductNode_Float66: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb7,SumNode_Float13Output_79,ProductNode_Float66Output_80);

ProductNode_Float67: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float67weight,v3,ProductNode_Float67Output_81);

ProductNode_Float68: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float68weight,ProductNode_Float4Output_5,ProductNode_Float68Output_82);

ProductNode_Float69: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float69weight,ProductNode_Float16Output_19,ProductNode_Float69Output_83);

ProductNode_Float70: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float70weight,vb3,ProductNode_Float70Output_84);

ProductNode_Float71: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float71weight,ProductNode_Float7Output_8,ProductNode_Float71Output_85);

ProductNode_Float72: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float72weight,ProductNode_Float19Output_22,ProductNode_Float72Output_86);

SumNode_Float14: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float72Output_86,ProductNode_Float69Output_83,SumNode_Float14Output_87);

ProductNode_Float73: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float14Output_87,ProductNode_Float66Output_80,ProductNode_Float73Output_88);

ProductNode_Float74: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float74weight,ProductNode_Float73Output_88,ProductNode_Float74Output_89);

SumNode_Float15: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float74Output_89,ProductNode_Float63Output_76,SumNode_Float15Output_90);

ProductNode_Float75: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float15Output_90,ProductNode_Float0Output_0,ProductNode_Float75Output_91);

ProductNode_Float76: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float76weight,ProductNode_Float75Output_91,ProductNode_Float76Output_92);

ProductNode_Float77: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float77weight,vb4,ProductNode_Float77Output_93);

ProductNode_Float78: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float78weight,v8,ProductNode_Float78Output_94);

ProductNode_Float79: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float79weight,vb8,ProductNode_Float79Output_95);

SumNode_Float16: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float79Output_95,ProductNode_Float78Output_94,SumNode_Float16Output_96);

ProductNode_Float80: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v7,SumNode_Float16Output_96,ProductNode_Float80Output_97);

ProductNode_Float81: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float81weight,v3,ProductNode_Float81Output_98);

ProductNode_Float82: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float82weight,ProductNode_Float29Output_35,ProductNode_Float82Output_99);

ProductNode_Float83: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float83weight,ProductNode_Float30Output_36,ProductNode_Float83Output_100);

ProductNode_Float84: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float84weight,vb3,ProductNode_Float84Output_101);

ProductNode_Float85: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float85weight,ProductNode_Float32Output_38,ProductNode_Float85Output_102);

ProductNode_Float86: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float86weight,ProductNode_Float33Output_39,ProductNode_Float86Output_103);

SumNode_Float17: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float86Output_103,ProductNode_Float83Output_100,SumNode_Float17Output_104);

ProductNode_Float87: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float17Output_104,ProductNode_Float80Output_97,ProductNode_Float87Output_105);

ProductNode_Float88: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float88weight,ProductNode_Float87Output_105,ProductNode_Float88Output_106);

ProductNode_Float89: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float89weight,v8,ProductNode_Float89Output_107);

ProductNode_Float90: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float90weight,vb8,ProductNode_Float90Output_108);

SumNode_Float18: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float90Output_108,ProductNode_Float89Output_107,SumNode_Float18Output_109);

ProductNode_Float91: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb7,SumNode_Float18Output_109,ProductNode_Float91Output_110);

ProductNode_Float92: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float92weight,v3,ProductNode_Float92Output_111);

ProductNode_Float93: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float93weight,ProductNode_Float29Output_35,ProductNode_Float93Output_112);

ProductNode_Float94: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float94weight,ProductNode_Float41Output_49,ProductNode_Float94Output_113);

ProductNode_Float95: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float95weight,vb3,ProductNode_Float95Output_114);

ProductNode_Float96: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float96weight,ProductNode_Float32Output_38,ProductNode_Float96Output_115);

ProductNode_Float97: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float97weight,ProductNode_Float44Output_52,ProductNode_Float97Output_116);

SumNode_Float19: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float97Output_116,ProductNode_Float94Output_113,SumNode_Float19Output_117);

ProductNode_Float98: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float19Output_117,ProductNode_Float91Output_110,ProductNode_Float98Output_118);

ProductNode_Float99: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float99weight,ProductNode_Float98Output_118,ProductNode_Float99Output_119);

SumNode_Float20: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float99Output_119,ProductNode_Float88Output_106,SumNode_Float20Output_120);

ProductNode_Float100: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float20Output_120,ProductNode_Float25Output_30,ProductNode_Float100Output_121);

ProductNode_Float101: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float101weight,ProductNode_Float100Output_121,ProductNode_Float101Output_122);

SumNode_Float21: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float101Output_122,ProductNode_Float76Output_92,SumNode_Float21Output_123);

ProductNode_Float102: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb5,SumNode_Float21Output_123,ProductNode_Float102Output_124);

ProductNode_Float103: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float103weight,ProductNode_Float102Output_124,ProductNode_Float103Output_125);

SumNode_Float22: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float103Output_125,ProductNode_Float51Output_62,SumNode_Float22Output_126);

ProductNode_Float104: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v16,SumNode_Float22Output_126,ProductNode_Float104Output_127);

ProductNode_Float105: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float105weight,v11,ProductNode_Float105Output_128);

ProductNode_Float106: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float106weight,vb11,ProductNode_Float106Output_129);

SumNode_Float23: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float106Output_129,ProductNode_Float105Output_128,SumNode_Float23Output_130);

ProductNode_Float107: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v12,SumNode_Float23Output_130,ProductNode_Float107Output_131);

ProductNode_Float108: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float108weight,ProductNode_Float107Output_131,ProductNode_Float108Output_132);

ProductNode_Float109: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float109weight,v2,ProductNode_Float109Output_133);

ProductNode_Float110: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float110weight,vb2,ProductNode_Float110Output_134);

SumNode_Float24: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float110Output_134,ProductNode_Float109Output_133,SumNode_Float24Output_135);

ProductNode_Float111: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float24Output_135,ProductNode_Float108Output_132,ProductNode_Float111Output_136);

ProductNode_Float112: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float112weight,v11,ProductNode_Float112Output_137);

ProductNode_Float113: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float113weight,vb11,ProductNode_Float113Output_138);

SumNode_Float25: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float113Output_138,ProductNode_Float112Output_137,SumNode_Float25Output_139);

ProductNode_Float114: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb12,SumNode_Float25Output_139,ProductNode_Float114Output_140);

ProductNode_Float115: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float115weight,ProductNode_Float114Output_140,ProductNode_Float115Output_141);

ProductNode_Float116: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float116weight,v2,ProductNode_Float116Output_142);

ProductNode_Float117: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float117weight,vb2,ProductNode_Float117Output_143);

SumNode_Float26: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float117Output_143,ProductNode_Float116Output_142,SumNode_Float26Output_144);

ProductNode_Float118: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float26Output_144,ProductNode_Float115Output_141,ProductNode_Float118Output_145);

SumNode_Float27: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float118Output_145,ProductNode_Float111Output_136,SumNode_Float27Output_146);

ProductNode_Float119: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v13,SumNode_Float27Output_146,ProductNode_Float119Output_147);

ProductNode_Float120: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float120weight,ProductNode_Float119Output_147,ProductNode_Float120Output_148);

ProductNode_Float121: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float121weight,v11,ProductNode_Float121Output_149);

ProductNode_Float122: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float122weight,vb11,ProductNode_Float122Output_150);

SumNode_Float28: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float122Output_150,ProductNode_Float121Output_149,SumNode_Float28Output_151);

ProductNode_Float123: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v12,SumNode_Float28Output_151,ProductNode_Float123Output_152);

ProductNode_Float124: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float124weight,ProductNode_Float123Output_152,ProductNode_Float124Output_153);

ProductNode_Float125: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float125weight,v2,ProductNode_Float125Output_154);

ProductNode_Float126: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float126weight,vb2,ProductNode_Float126Output_155);

SumNode_Float29: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float126Output_155,ProductNode_Float125Output_154,SumNode_Float29Output_156);

ProductNode_Float127: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float29Output_156,ProductNode_Float124Output_153,ProductNode_Float127Output_157);

ProductNode_Float128: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float128weight,v11,ProductNode_Float128Output_158);

ProductNode_Float129: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float129weight,vb11,ProductNode_Float129Output_159);

SumNode_Float30: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float129Output_159,ProductNode_Float128Output_158,SumNode_Float30Output_160);

ProductNode_Float130: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb12,SumNode_Float30Output_160,ProductNode_Float130Output_161);

ProductNode_Float131: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float131weight,ProductNode_Float130Output_161,ProductNode_Float131Output_162);

ProductNode_Float132: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float132weight,v2,ProductNode_Float132Output_163);

ProductNode_Float133: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float133weight,vb2,ProductNode_Float133Output_164);

SumNode_Float31: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float133Output_164,ProductNode_Float132Output_163,SumNode_Float31Output_165);

ProductNode_Float134: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float31Output_165,ProductNode_Float131Output_162,ProductNode_Float134Output_166);

SumNode_Float32: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float134Output_166,ProductNode_Float127Output_157,SumNode_Float32Output_167);

ProductNode_Float135: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb13,SumNode_Float32Output_167,ProductNode_Float135Output_168);

ProductNode_Float136: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float136weight,ProductNode_Float135Output_168,ProductNode_Float136Output_169);

SumNode_Float33: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float136Output_169,ProductNode_Float120Output_148,SumNode_Float33Output_170);

ProductNode_Float137: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v10,SumNode_Float33Output_170,ProductNode_Float137Output_171);

ProductNode_Float138: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float138weight,v1,ProductNode_Float138Output_172);

ProductNode_Float139: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float139weight,vb1,ProductNode_Float139Output_173);

SumNode_Float34: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float139Output_173,ProductNode_Float138Output_172,SumNode_Float34Output_174);

ProductNode_Float140: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v9,SumNode_Float34Output_174,ProductNode_Float140Output_175);

ProductNode_Float141: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float141weight,ProductNode_Float140Output_175,ProductNode_Float141Output_176);

ProductNode_Float142: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float142weight,ProductNode_Float141Output_176,ProductNode_Float142Output_177);

ProductNode_Float143: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float143weight,v1,ProductNode_Float143Output_178);

ProductNode_Float144: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float144weight,vb1,ProductNode_Float144Output_179);

SumNode_Float35: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float144Output_179,ProductNode_Float143Output_178,SumNode_Float35Output_180);

ProductNode_Float145: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb9,SumNode_Float35Output_180,ProductNode_Float145Output_181);

ProductNode_Float146: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float146weight,ProductNode_Float145Output_181,ProductNode_Float146Output_182);

ProductNode_Float147: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float147weight,ProductNode_Float146Output_182,ProductNode_Float147Output_183);

SumNode_Float36: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float147Output_183,ProductNode_Float142Output_177,SumNode_Float36Output_184);

ProductNode_Float148: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float36Output_184,ProductNode_Float137Output_171,ProductNode_Float148Output_185);

ProductNode_Float149: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float149weight,v11,ProductNode_Float149Output_186);

ProductNode_Float150: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float150weight,vb11,ProductNode_Float150Output_187);

SumNode_Float37: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float106Output_129,ProductNode_Float105Output_128,SumNode_Float37Output_188);

ProductNode_Float151: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v12,SumNode_Float23Output_130,ProductNode_Float151Output_189);

ProductNode_Float152: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float152weight,ProductNode_Float107Output_131,ProductNode_Float152Output_190);

ProductNode_Float153: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float153weight,v2,ProductNode_Float153Output_191);

ProductNode_Float154: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float154weight,vb2,ProductNode_Float154Output_192);

SumNode_Float38: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float110Output_134,ProductNode_Float109Output_133,SumNode_Float38Output_193);

ProductNode_Float155: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float24Output_135,ProductNode_Float108Output_132,ProductNode_Float155Output_194);

ProductNode_Float156: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float156weight,v11,ProductNode_Float156Output_195);

ProductNode_Float157: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float157weight,vb11,ProductNode_Float157Output_196);

SumNode_Float39: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float113Output_138,ProductNode_Float112Output_137,SumNode_Float39Output_197);

ProductNode_Float158: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb12,SumNode_Float25Output_139,ProductNode_Float158Output_198);

ProductNode_Float159: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float159weight,ProductNode_Float114Output_140,ProductNode_Float159Output_199);

ProductNode_Float160: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float160weight,v2,ProductNode_Float160Output_200);

ProductNode_Float161: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float161weight,vb2,ProductNode_Float161Output_201);

SumNode_Float40: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float117Output_143,ProductNode_Float116Output_142,SumNode_Float40Output_202);

ProductNode_Float162: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float26Output_144,ProductNode_Float115Output_141,ProductNode_Float162Output_203);

SumNode_Float41: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float118Output_145,ProductNode_Float111Output_136,SumNode_Float41Output_204);

ProductNode_Float163: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v13,SumNode_Float27Output_146,ProductNode_Float163Output_205);

ProductNode_Float164: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float164weight,ProductNode_Float119Output_147,ProductNode_Float164Output_206);

ProductNode_Float165: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float165weight,v11,ProductNode_Float165Output_207);

ProductNode_Float166: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float166weight,vb11,ProductNode_Float166Output_208);

SumNode_Float42: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float122Output_150,ProductNode_Float121Output_149,SumNode_Float42Output_209);

ProductNode_Float167: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v12,SumNode_Float28Output_151,ProductNode_Float167Output_210);

ProductNode_Float168: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float168weight,ProductNode_Float123Output_152,ProductNode_Float168Output_211);

ProductNode_Float169: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float169weight,v2,ProductNode_Float169Output_212);

ProductNode_Float170: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float170weight,vb2,ProductNode_Float170Output_213);

SumNode_Float43: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float126Output_155,ProductNode_Float125Output_154,SumNode_Float43Output_214);

ProductNode_Float171: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float29Output_156,ProductNode_Float124Output_153,ProductNode_Float171Output_215);

ProductNode_Float172: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float172weight,v11,ProductNode_Float172Output_216);

ProductNode_Float173: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float173weight,vb11,ProductNode_Float173Output_217);

SumNode_Float44: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float129Output_159,ProductNode_Float128Output_158,SumNode_Float44Output_218);

ProductNode_Float174: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb12,SumNode_Float30Output_160,ProductNode_Float174Output_219);

ProductNode_Float175: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float175weight,ProductNode_Float130Output_161,ProductNode_Float175Output_220);

ProductNode_Float176: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float176weight,v2,ProductNode_Float176Output_221);

ProductNode_Float177: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float177weight,vb2,ProductNode_Float177Output_222);

SumNode_Float45: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float133Output_164,ProductNode_Float132Output_163,SumNode_Float45Output_223);

ProductNode_Float178: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float31Output_165,ProductNode_Float131Output_162,ProductNode_Float178Output_224);

SumNode_Float46: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float134Output_166,ProductNode_Float127Output_157,SumNode_Float46Output_225);

ProductNode_Float179: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb13,SumNode_Float32Output_167,ProductNode_Float179Output_226);

ProductNode_Float180: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float180weight,ProductNode_Float135Output_168,ProductNode_Float180Output_227);

SumNode_Float47: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float180Output_227,ProductNode_Float164Output_206,SumNode_Float47Output_228);

ProductNode_Float181: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb10,SumNode_Float47Output_228,ProductNode_Float181Output_229);

ProductNode_Float182: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float182weight,v1,ProductNode_Float182Output_230);

ProductNode_Float183: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float183weight,vb1,ProductNode_Float183Output_231);

SumNode_Float48: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float183Output_231,ProductNode_Float182Output_230,SumNode_Float48Output_232);

ProductNode_Float184: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v9,SumNode_Float48Output_232,ProductNode_Float184Output_233);

ProductNode_Float185: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float185weight,ProductNode_Float184Output_233,ProductNode_Float185Output_234);

ProductNode_Float186: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float186weight,ProductNode_Float185Output_234,ProductNode_Float186Output_235);

ProductNode_Float187: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float187weight,v1,ProductNode_Float187Output_236);

ProductNode_Float188: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float188weight,vb1,ProductNode_Float188Output_237);

SumNode_Float49: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float188Output_237,ProductNode_Float187Output_236,SumNode_Float49Output_238);

ProductNode_Float189: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb9,SumNode_Float49Output_238,ProductNode_Float189Output_239);

ProductNode_Float190: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float190weight,ProductNode_Float189Output_239,ProductNode_Float190Output_240);

ProductNode_Float191: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float191weight,ProductNode_Float190Output_240,ProductNode_Float191Output_241);

SumNode_Float50: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float191Output_241,ProductNode_Float186Output_235,SumNode_Float50Output_242);

ProductNode_Float192: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float50Output_242,ProductNode_Float181Output_229,ProductNode_Float192Output_243);

SumNode_Float51: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float192Output_243,ProductNode_Float148Output_185,SumNode_Float51Output_244);

ProductNode_Float193: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v15,SumNode_Float51Output_244,ProductNode_Float193Output_245);

ProductNode_Float194: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float194weight,ProductNode_Float193Output_245,ProductNode_Float194Output_246);

ProductNode_Float195: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float195weight,v11,ProductNode_Float195Output_247);

ProductNode_Float196: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float196weight,vb11,ProductNode_Float196Output_248);

SumNode_Float52: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float106Output_129,ProductNode_Float105Output_128,SumNode_Float52Output_249);

ProductNode_Float197: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v12,SumNode_Float23Output_130,ProductNode_Float197Output_250);

ProductNode_Float198: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float198weight,ProductNode_Float107Output_131,ProductNode_Float198Output_251);

ProductNode_Float199: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float199weight,v2,ProductNode_Float199Output_252);

ProductNode_Float200: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float200weight,vb2,ProductNode_Float200Output_253);

SumNode_Float53: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float200Output_253,ProductNode_Float199Output_252,SumNode_Float53Output_254);

ProductNode_Float201: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float53Output_254,ProductNode_Float108Output_132,ProductNode_Float201Output_255);

ProductNode_Float202: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float202weight,v11,ProductNode_Float202Output_256);

ProductNode_Float203: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float203weight,vb11,ProductNode_Float203Output_257);

SumNode_Float54: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float113Output_138,ProductNode_Float112Output_137,SumNode_Float54Output_258);

ProductNode_Float204: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb12,SumNode_Float25Output_139,ProductNode_Float204Output_259);

ProductNode_Float205: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float205weight,ProductNode_Float114Output_140,ProductNode_Float205Output_260);

ProductNode_Float206: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float206weight,v2,ProductNode_Float206Output_261);

ProductNode_Float207: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float207weight,vb2,ProductNode_Float207Output_262);

SumNode_Float55: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float207Output_262,ProductNode_Float206Output_261,SumNode_Float55Output_263);

ProductNode_Float208: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float55Output_263,ProductNode_Float115Output_141,ProductNode_Float208Output_264);

SumNode_Float56: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float208Output_264,ProductNode_Float201Output_255,SumNode_Float56Output_265);

ProductNode_Float209: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v13,SumNode_Float56Output_265,ProductNode_Float209Output_266);

ProductNode_Float210: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float210weight,ProductNode_Float209Output_266,ProductNode_Float210Output_267);

ProductNode_Float211: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float211weight,v11,ProductNode_Float211Output_268);

ProductNode_Float212: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float212weight,vb11,ProductNode_Float212Output_269);

SumNode_Float57: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float122Output_150,ProductNode_Float121Output_149,SumNode_Float57Output_270);

ProductNode_Float213: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v12,SumNode_Float28Output_151,ProductNode_Float213Output_271);

ProductNode_Float214: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float214weight,ProductNode_Float123Output_152,ProductNode_Float214Output_272);

ProductNode_Float215: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float215weight,v2,ProductNode_Float215Output_273);

ProductNode_Float216: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float216weight,vb2,ProductNode_Float216Output_274);

SumNode_Float58: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float216Output_274,ProductNode_Float215Output_273,SumNode_Float58Output_275);

ProductNode_Float217: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float58Output_275,ProductNode_Float124Output_153,ProductNode_Float217Output_276);

ProductNode_Float218: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float218weight,v11,ProductNode_Float218Output_277);

ProductNode_Float219: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float219weight,vb11,ProductNode_Float219Output_278);

SumNode_Float59: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float129Output_159,ProductNode_Float128Output_158,SumNode_Float59Output_279);

ProductNode_Float220: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb12,SumNode_Float30Output_160,ProductNode_Float220Output_280);

ProductNode_Float221: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float221weight,ProductNode_Float130Output_161,ProductNode_Float221Output_281);

ProductNode_Float222: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float222weight,v2,ProductNode_Float222Output_282);

ProductNode_Float223: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float223weight,vb2,ProductNode_Float223Output_283);

SumNode_Float60: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float223Output_283,ProductNode_Float222Output_282,SumNode_Float60Output_284);

ProductNode_Float224: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float60Output_284,ProductNode_Float131Output_162,ProductNode_Float224Output_285);

SumNode_Float61: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float224Output_285,ProductNode_Float217Output_276,SumNode_Float61Output_286);

ProductNode_Float225: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb13,SumNode_Float61Output_286,ProductNode_Float225Output_287);

ProductNode_Float226: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float226weight,ProductNode_Float225Output_287,ProductNode_Float226Output_288);

SumNode_Float62: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float226Output_288,ProductNode_Float210Output_267,SumNode_Float62Output_289);

ProductNode_Float227: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v10,SumNode_Float62Output_289,ProductNode_Float227Output_290);

ProductNode_Float228: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float228weight,v1,ProductNode_Float228Output_291);

ProductNode_Float229: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float229weight,vb1,ProductNode_Float229Output_292);

SumNode_Float63: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float139Output_173,ProductNode_Float138Output_172,SumNode_Float63Output_293);

ProductNode_Float230: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v9,SumNode_Float34Output_174,ProductNode_Float230Output_294);

ProductNode_Float231: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float231weight,ProductNode_Float140Output_175,ProductNode_Float231Output_295);

ProductNode_Float232: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float232weight,ProductNode_Float231Output_295,ProductNode_Float232Output_296);

ProductNode_Float233: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float233weight,v1,ProductNode_Float233Output_297);

ProductNode_Float234: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float234weight,vb1,ProductNode_Float234Output_298);

SumNode_Float64: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float144Output_179,ProductNode_Float143Output_178,SumNode_Float64Output_299);

ProductNode_Float235: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb9,SumNode_Float35Output_180,ProductNode_Float235Output_300);

ProductNode_Float236: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float236weight,ProductNode_Float145Output_181,ProductNode_Float236Output_301);

ProductNode_Float237: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float237weight,ProductNode_Float236Output_301,ProductNode_Float237Output_302);

SumNode_Float65: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float237Output_302,ProductNode_Float232Output_296,SumNode_Float65Output_303);

ProductNode_Float238: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float65Output_303,ProductNode_Float227Output_290,ProductNode_Float238Output_304);

ProductNode_Float239: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float239weight,v11,ProductNode_Float239Output_305);

ProductNode_Float240: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float240weight,vb11,ProductNode_Float240Output_306);

SumNode_Float66: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float106Output_129,ProductNode_Float105Output_128,SumNode_Float66Output_307);

ProductNode_Float241: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v12,SumNode_Float23Output_130,ProductNode_Float241Output_308);

ProductNode_Float242: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float242weight,ProductNode_Float107Output_131,ProductNode_Float242Output_309);

ProductNode_Float243: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float243weight,v2,ProductNode_Float243Output_310);

ProductNode_Float244: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float244weight,vb2,ProductNode_Float244Output_311);

SumNode_Float67: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float200Output_253,ProductNode_Float199Output_252,SumNode_Float67Output_312);

ProductNode_Float245: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float53Output_254,ProductNode_Float108Output_132,ProductNode_Float245Output_313);

ProductNode_Float246: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float246weight,v11,ProductNode_Float246Output_314);

ProductNode_Float247: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float247weight,vb11,ProductNode_Float247Output_315);

SumNode_Float68: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float113Output_138,ProductNode_Float112Output_137,SumNode_Float68Output_316);

ProductNode_Float248: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb12,SumNode_Float25Output_139,ProductNode_Float248Output_317);

ProductNode_Float249: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float249weight,ProductNode_Float114Output_140,ProductNode_Float249Output_318);

ProductNode_Float250: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float250weight,v2,ProductNode_Float250Output_319);

ProductNode_Float251: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float251weight,vb2,ProductNode_Float251Output_320);

SumNode_Float69: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float207Output_262,ProductNode_Float206Output_261,SumNode_Float69Output_321);

ProductNode_Float252: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float55Output_263,ProductNode_Float115Output_141,ProductNode_Float252Output_322);

SumNode_Float70: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float208Output_264,ProductNode_Float201Output_255,SumNode_Float70Output_323);

ProductNode_Float253: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v13,SumNode_Float56Output_265,ProductNode_Float253Output_324);

ProductNode_Float254: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float254weight,ProductNode_Float209Output_266,ProductNode_Float254Output_325);

ProductNode_Float255: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float255weight,v11,ProductNode_Float255Output_326);

ProductNode_Float256: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float256weight,vb11,ProductNode_Float256Output_327);

SumNode_Float71: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float122Output_150,ProductNode_Float121Output_149,SumNode_Float71Output_328);

ProductNode_Float257: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v12,SumNode_Float28Output_151,ProductNode_Float257Output_329);

ProductNode_Float258: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float258weight,ProductNode_Float123Output_152,ProductNode_Float258Output_330);

ProductNode_Float259: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float259weight,v2,ProductNode_Float259Output_331);

ProductNode_Float260: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float260weight,vb2,ProductNode_Float260Output_332);

SumNode_Float72: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float216Output_274,ProductNode_Float215Output_273,SumNode_Float72Output_333);

ProductNode_Float261: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float58Output_275,ProductNode_Float124Output_153,ProductNode_Float261Output_334);

ProductNode_Float262: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float262weight,v11,ProductNode_Float262Output_335);

ProductNode_Float263: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float263weight,vb11,ProductNode_Float263Output_336);

SumNode_Float73: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float129Output_159,ProductNode_Float128Output_158,SumNode_Float73Output_337);

ProductNode_Float264: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb12,SumNode_Float30Output_160,ProductNode_Float264Output_338);

ProductNode_Float265: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float265weight,ProductNode_Float130Output_161,ProductNode_Float265Output_339);

ProductNode_Float266: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float266weight,v2,ProductNode_Float266Output_340);

ProductNode_Float267: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float267weight,vb2,ProductNode_Float267Output_341);

SumNode_Float74: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float223Output_283,ProductNode_Float222Output_282,SumNode_Float74Output_342);

ProductNode_Float268: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float60Output_284,ProductNode_Float131Output_162,ProductNode_Float268Output_343);

SumNode_Float75: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float224Output_285,ProductNode_Float217Output_276,SumNode_Float75Output_344);

ProductNode_Float269: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb13,SumNode_Float61Output_286,ProductNode_Float269Output_345);

ProductNode_Float270: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float270weight,ProductNode_Float225Output_287,ProductNode_Float270Output_346);

SumNode_Float76: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float270Output_346,ProductNode_Float254Output_325,SumNode_Float76Output_347);

ProductNode_Float271: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb10,SumNode_Float76Output_347,ProductNode_Float271Output_348);

ProductNode_Float272: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float272weight,v1,ProductNode_Float272Output_349);

ProductNode_Float273: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float273weight,vb1,ProductNode_Float273Output_350);

SumNode_Float77: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float183Output_231,ProductNode_Float182Output_230,SumNode_Float77Output_351);

ProductNode_Float274: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v9,SumNode_Float48Output_232,ProductNode_Float274Output_352);

ProductNode_Float275: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float275weight,ProductNode_Float184Output_233,ProductNode_Float275Output_353);

ProductNode_Float276: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float276weight,ProductNode_Float275Output_353,ProductNode_Float276Output_354);

ProductNode_Float277: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float277weight,v1,ProductNode_Float277Output_355);

ProductNode_Float278: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float278weight,vb1,ProductNode_Float278Output_356);

SumNode_Float78: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float188Output_237,ProductNode_Float187Output_236,SumNode_Float78Output_357);

ProductNode_Float279: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb9,SumNode_Float49Output_238,ProductNode_Float279Output_358);

ProductNode_Float280: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float280weight,ProductNode_Float189Output_239,ProductNode_Float280Output_359);

ProductNode_Float281: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float281weight,ProductNode_Float280Output_359,ProductNode_Float281Output_360);

SumNode_Float79: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float281Output_360,ProductNode_Float276Output_354,SumNode_Float79Output_361);

ProductNode_Float282: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float79Output_361,ProductNode_Float271Output_348,ProductNode_Float282Output_362);

SumNode_Float80: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float282Output_362,ProductNode_Float238Output_304,SumNode_Float80Output_363);

ProductNode_Float283: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb15,SumNode_Float80Output_363,ProductNode_Float283Output_364);

ProductNode_Float284: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float284weight,ProductNode_Float283Output_364,ProductNode_Float284Output_365);

SumNode_Float81: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float284Output_365,ProductNode_Float194Output_246,SumNode_Float81Output_366);

ProductNode_Float285: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float81Output_366,ProductNode_Float104Output_127,ProductNode_Float285Output_367);

ProductNode_Float286: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float286weight,v4,ProductNode_Float286Output_368);

ProductNode_Float287: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float287weight,v8,ProductNode_Float287Output_369);

ProductNode_Float288: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float288weight,vb8,ProductNode_Float288Output_370);

SumNode_Float82: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2Output_2,ProductNode_Float1Output_1,SumNode_Float82Output_371);

ProductNode_Float289: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v7,SumNode_Float0Output_3,ProductNode_Float289Output_372);

ProductNode_Float290: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float290weight,v3,ProductNode_Float290Output_373);

ProductNode_Float291: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float291weight,ProductNode_Float4Output_5,ProductNode_Float291Output_374);

ProductNode_Float292: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float292weight,ProductNode_Float5Output_6,ProductNode_Float292Output_375);

ProductNode_Float293: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float293weight,vb3,ProductNode_Float293Output_376);

ProductNode_Float294: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float294weight,ProductNode_Float7Output_8,ProductNode_Float294Output_377);

ProductNode_Float295: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float295weight,ProductNode_Float8Output_9,ProductNode_Float295Output_378);

SumNode_Float83: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float9Output_10,ProductNode_Float6Output_7,SumNode_Float83Output_379);

ProductNode_Float296: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float1Output_11,ProductNode_Float3Output_4,ProductNode_Float296Output_380);

ProductNode_Float297: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float297weight,ProductNode_Float10Output_12,ProductNode_Float297Output_381);

ProductNode_Float298: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float298weight,v8,ProductNode_Float298Output_382);

ProductNode_Float299: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float299weight,vb8,ProductNode_Float299Output_383);

SumNode_Float84: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float13Output_15,ProductNode_Float12Output_14,SumNode_Float84Output_384);

ProductNode_Float300: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb7,SumNode_Float2Output_16,ProductNode_Float300Output_385);

ProductNode_Float301: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float301weight,v3,ProductNode_Float301Output_386);

ProductNode_Float302: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float302weight,ProductNode_Float4Output_5,ProductNode_Float302Output_387);

ProductNode_Float303: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float303weight,ProductNode_Float16Output_19,ProductNode_Float303Output_388);

ProductNode_Float304: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float304weight,vb3,ProductNode_Float304Output_389);

ProductNode_Float305: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float305weight,ProductNode_Float7Output_8,ProductNode_Float305Output_390);

ProductNode_Float306: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float306weight,ProductNode_Float19Output_22,ProductNode_Float306Output_391);

SumNode_Float85: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float20Output_23,ProductNode_Float17Output_20,SumNode_Float85Output_392);

ProductNode_Float307: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float3Output_24,ProductNode_Float14Output_17,ProductNode_Float307Output_393);

ProductNode_Float308: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float308weight,ProductNode_Float21Output_25,ProductNode_Float308Output_394);

SumNode_Float86: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float22Output_26,ProductNode_Float11Output_13,SumNode_Float86Output_395);

ProductNode_Float309: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float4Output_27,ProductNode_Float0Output_0,ProductNode_Float309Output_396);

ProductNode_Float310: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float310weight,ProductNode_Float23Output_28,ProductNode_Float310Output_397);

ProductNode_Float311: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float311weight,vb4,ProductNode_Float311Output_398);

ProductNode_Float312: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float312weight,v8,ProductNode_Float312Output_399);

ProductNode_Float313: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float313weight,vb8,ProductNode_Float313Output_400);

SumNode_Float87: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float27Output_32,ProductNode_Float26Output_31,SumNode_Float87Output_401);

ProductNode_Float314: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v7,SumNode_Float5Output_33,ProductNode_Float314Output_402);

ProductNode_Float315: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float315weight,v3,ProductNode_Float315Output_403);

ProductNode_Float316: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float316weight,ProductNode_Float29Output_35,ProductNode_Float316Output_404);

ProductNode_Float317: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float317weight,ProductNode_Float30Output_36,ProductNode_Float317Output_405);

ProductNode_Float318: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float318weight,vb3,ProductNode_Float318Output_406);

ProductNode_Float319: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float319weight,ProductNode_Float32Output_38,ProductNode_Float319Output_407);

ProductNode_Float320: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float320weight,ProductNode_Float33Output_39,ProductNode_Float320Output_408);

SumNode_Float88: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float34Output_40,ProductNode_Float31Output_37,SumNode_Float88Output_409);

ProductNode_Float321: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float6Output_41,ProductNode_Float28Output_34,ProductNode_Float321Output_410);

ProductNode_Float322: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float322weight,ProductNode_Float35Output_42,ProductNode_Float322Output_411);

ProductNode_Float323: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float323weight,v8,ProductNode_Float323Output_412);

ProductNode_Float324: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float324weight,vb8,ProductNode_Float324Output_413);

SumNode_Float89: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float38Output_45,ProductNode_Float37Output_44,SumNode_Float89Output_414);

ProductNode_Float325: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb7,SumNode_Float7Output_46,ProductNode_Float325Output_415);

ProductNode_Float326: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float326weight,v3,ProductNode_Float326Output_416);

ProductNode_Float327: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float327weight,ProductNode_Float29Output_35,ProductNode_Float327Output_417);

ProductNode_Float328: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float328weight,ProductNode_Float41Output_49,ProductNode_Float328Output_418);

ProductNode_Float329: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float329weight,vb3,ProductNode_Float329Output_419);

ProductNode_Float330: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float330weight,ProductNode_Float32Output_38,ProductNode_Float330Output_420);

ProductNode_Float331: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float331weight,ProductNode_Float44Output_52,ProductNode_Float331Output_421);

SumNode_Float90: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float45Output_53,ProductNode_Float42Output_50,SumNode_Float90Output_422);

ProductNode_Float332: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float8Output_54,ProductNode_Float39Output_47,ProductNode_Float332Output_423);

ProductNode_Float333: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float333weight,ProductNode_Float46Output_55,ProductNode_Float333Output_424);

SumNode_Float91: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float47Output_56,ProductNode_Float36Output_43,SumNode_Float91Output_425);

ProductNode_Float334: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float9Output_57,ProductNode_Float25Output_30,ProductNode_Float334Output_426);

ProductNode_Float335: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float335weight,ProductNode_Float48Output_58,ProductNode_Float335Output_427);

SumNode_Float92: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float335Output_427,ProductNode_Float310Output_397,SumNode_Float92Output_428);

ProductNode_Float336: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v5,SumNode_Float92Output_428,ProductNode_Float336Output_429);

ProductNode_Float337: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float337weight,ProductNode_Float336Output_429,ProductNode_Float337Output_430);

ProductNode_Float338: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float338weight,v4,ProductNode_Float338Output_431);

ProductNode_Float339: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float339weight,v8,ProductNode_Float339Output_432);

ProductNode_Float340: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float340weight,vb8,ProductNode_Float340Output_433);

SumNode_Float93: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float54Output_65,ProductNode_Float53Output_64,SumNode_Float93Output_434);

ProductNode_Float341: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v7,SumNode_Float11Output_66,ProductNode_Float341Output_435);

ProductNode_Float342: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float342weight,v3,ProductNode_Float342Output_436);

ProductNode_Float343: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float343weight,ProductNode_Float4Output_5,ProductNode_Float343Output_437);

ProductNode_Float344: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float344weight,ProductNode_Float5Output_6,ProductNode_Float344Output_438);

ProductNode_Float345: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float345weight,vb3,ProductNode_Float345Output_439);

ProductNode_Float346: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float346weight,ProductNode_Float7Output_8,ProductNode_Float346Output_440);

ProductNode_Float347: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float347weight,ProductNode_Float8Output_9,ProductNode_Float347Output_441);

SumNode_Float94: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float61Output_73,ProductNode_Float58Output_70,SumNode_Float94Output_442);

ProductNode_Float348: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float12Output_74,ProductNode_Float55Output_67,ProductNode_Float348Output_443);

ProductNode_Float349: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float349weight,ProductNode_Float62Output_75,ProductNode_Float349Output_444);

ProductNode_Float350: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float350weight,v8,ProductNode_Float350Output_445);

ProductNode_Float351: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float351weight,vb8,ProductNode_Float351Output_446);

SumNode_Float95: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float65Output_78,ProductNode_Float64Output_77,SumNode_Float95Output_447);

ProductNode_Float352: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb7,SumNode_Float13Output_79,ProductNode_Float352Output_448);

ProductNode_Float353: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float353weight,v3,ProductNode_Float353Output_449);

ProductNode_Float354: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float354weight,ProductNode_Float4Output_5,ProductNode_Float354Output_450);

ProductNode_Float355: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float355weight,ProductNode_Float16Output_19,ProductNode_Float355Output_451);

ProductNode_Float356: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float356weight,vb3,ProductNode_Float356Output_452);

ProductNode_Float357: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float357weight,ProductNode_Float7Output_8,ProductNode_Float357Output_453);

ProductNode_Float358: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float358weight,ProductNode_Float19Output_22,ProductNode_Float358Output_454);

SumNode_Float96: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float72Output_86,ProductNode_Float69Output_83,SumNode_Float96Output_455);

ProductNode_Float359: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float14Output_87,ProductNode_Float66Output_80,ProductNode_Float359Output_456);

ProductNode_Float360: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float360weight,ProductNode_Float73Output_88,ProductNode_Float360Output_457);

SumNode_Float97: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float74Output_89,ProductNode_Float63Output_76,SumNode_Float97Output_458);

ProductNode_Float361: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float15Output_90,ProductNode_Float0Output_0,ProductNode_Float361Output_459);

ProductNode_Float362: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float362weight,ProductNode_Float75Output_91,ProductNode_Float362Output_460);

ProductNode_Float363: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float363weight,vb4,ProductNode_Float363Output_461);

ProductNode_Float364: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float364weight,v8,ProductNode_Float364Output_462);

ProductNode_Float365: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float365weight,vb8,ProductNode_Float365Output_463);

SumNode_Float98: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float79Output_95,ProductNode_Float78Output_94,SumNode_Float98Output_464);

ProductNode_Float366: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v7,SumNode_Float16Output_96,ProductNode_Float366Output_465);

ProductNode_Float367: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float367weight,v3,ProductNode_Float367Output_466);

ProductNode_Float368: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float368weight,ProductNode_Float29Output_35,ProductNode_Float368Output_467);

ProductNode_Float369: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float369weight,ProductNode_Float30Output_36,ProductNode_Float369Output_468);

ProductNode_Float370: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float370weight,vb3,ProductNode_Float370Output_469);

ProductNode_Float371: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float371weight,ProductNode_Float32Output_38,ProductNode_Float371Output_470);

ProductNode_Float372: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float372weight,ProductNode_Float33Output_39,ProductNode_Float372Output_471);

SumNode_Float99: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float86Output_103,ProductNode_Float83Output_100,SumNode_Float99Output_472);

ProductNode_Float373: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float17Output_104,ProductNode_Float80Output_97,ProductNode_Float373Output_473);

ProductNode_Float374: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float374weight,ProductNode_Float87Output_105,ProductNode_Float374Output_474);

ProductNode_Float375: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float375weight,v8,ProductNode_Float375Output_475);

ProductNode_Float376: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float376weight,vb8,ProductNode_Float376Output_476);

SumNode_Float100: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float90Output_108,ProductNode_Float89Output_107,SumNode_Float100Output_477);

ProductNode_Float377: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb7,SumNode_Float18Output_109,ProductNode_Float377Output_478);

ProductNode_Float378: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float378weight,v3,ProductNode_Float378Output_479);

ProductNode_Float379: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float379weight,ProductNode_Float29Output_35,ProductNode_Float379Output_480);

ProductNode_Float380: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float380weight,ProductNode_Float41Output_49,ProductNode_Float380Output_481);

ProductNode_Float381: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float381weight,vb3,ProductNode_Float381Output_482);

ProductNode_Float382: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float382weight,ProductNode_Float32Output_38,ProductNode_Float382Output_483);

ProductNode_Float383: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float383weight,ProductNode_Float44Output_52,ProductNode_Float383Output_484);

SumNode_Float101: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float97Output_116,ProductNode_Float94Output_113,SumNode_Float101Output_485);

ProductNode_Float384: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float19Output_117,ProductNode_Float91Output_110,ProductNode_Float384Output_486);

ProductNode_Float385: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float385weight,ProductNode_Float98Output_118,ProductNode_Float385Output_487);

SumNode_Float102: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float99Output_119,ProductNode_Float88Output_106,SumNode_Float102Output_488);

ProductNode_Float386: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float20Output_120,ProductNode_Float25Output_30,ProductNode_Float386Output_489);

ProductNode_Float387: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float387weight,ProductNode_Float100Output_121,ProductNode_Float387Output_490);

SumNode_Float103: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float387Output_490,ProductNode_Float362Output_460,SumNode_Float103Output_491);

ProductNode_Float388: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb5,SumNode_Float103Output_491,ProductNode_Float388Output_492);

ProductNode_Float389: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float389weight,ProductNode_Float388Output_492,ProductNode_Float389Output_493);

SumNode_Float104: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float389Output_493,ProductNode_Float337Output_430,SumNode_Float104Output_494);

ProductNode_Float390: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb16,SumNode_Float104Output_494,ProductNode_Float390Output_495);

ProductNode_Float391: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float391weight,v11,ProductNode_Float391Output_496);

ProductNode_Float392: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float392weight,vb11,ProductNode_Float392Output_497);

SumNode_Float105: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float106Output_129,ProductNode_Float105Output_128,SumNode_Float105Output_498);

ProductNode_Float393: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v12,SumNode_Float23Output_130,ProductNode_Float393Output_499);

ProductNode_Float394: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float394weight,ProductNode_Float107Output_131,ProductNode_Float394Output_500);

ProductNode_Float395: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float395weight,v2,ProductNode_Float395Output_501);

ProductNode_Float396: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float396weight,vb2,ProductNode_Float396Output_502);

SumNode_Float106: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float110Output_134,ProductNode_Float109Output_133,SumNode_Float106Output_503);

ProductNode_Float397: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float24Output_135,ProductNode_Float108Output_132,ProductNode_Float397Output_504);

ProductNode_Float398: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float398weight,v11,ProductNode_Float398Output_505);

ProductNode_Float399: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float399weight,vb11,ProductNode_Float399Output_506);

SumNode_Float107: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float113Output_138,ProductNode_Float112Output_137,SumNode_Float107Output_507);

ProductNode_Float400: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb12,SumNode_Float25Output_139,ProductNode_Float400Output_508);

ProductNode_Float401: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float401weight,ProductNode_Float114Output_140,ProductNode_Float401Output_509);

ProductNode_Float402: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float402weight,v2,ProductNode_Float402Output_510);

ProductNode_Float403: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float403weight,vb2,ProductNode_Float403Output_511);

SumNode_Float108: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float117Output_143,ProductNode_Float116Output_142,SumNode_Float108Output_512);

ProductNode_Float404: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float26Output_144,ProductNode_Float115Output_141,ProductNode_Float404Output_513);

SumNode_Float109: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float118Output_145,ProductNode_Float111Output_136,SumNode_Float109Output_514);

ProductNode_Float405: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v13,SumNode_Float27Output_146,ProductNode_Float405Output_515);

ProductNode_Float406: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float406weight,ProductNode_Float119Output_147,ProductNode_Float406Output_516);

ProductNode_Float407: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float407weight,v11,ProductNode_Float407Output_517);

ProductNode_Float408: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float408weight,vb11,ProductNode_Float408Output_518);

SumNode_Float110: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float122Output_150,ProductNode_Float121Output_149,SumNode_Float110Output_519);

ProductNode_Float409: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v12,SumNode_Float28Output_151,ProductNode_Float409Output_520);

ProductNode_Float410: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float410weight,ProductNode_Float123Output_152,ProductNode_Float410Output_521);

ProductNode_Float411: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float411weight,v2,ProductNode_Float411Output_522);

ProductNode_Float412: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float412weight,vb2,ProductNode_Float412Output_523);

SumNode_Float111: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float126Output_155,ProductNode_Float125Output_154,SumNode_Float111Output_524);

ProductNode_Float413: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float29Output_156,ProductNode_Float124Output_153,ProductNode_Float413Output_525);

ProductNode_Float414: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float414weight,v11,ProductNode_Float414Output_526);

ProductNode_Float415: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float415weight,vb11,ProductNode_Float415Output_527);

SumNode_Float112: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float129Output_159,ProductNode_Float128Output_158,SumNode_Float112Output_528);

ProductNode_Float416: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb12,SumNode_Float30Output_160,ProductNode_Float416Output_529);

ProductNode_Float417: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float417weight,ProductNode_Float130Output_161,ProductNode_Float417Output_530);

ProductNode_Float418: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float418weight,v2,ProductNode_Float418Output_531);

ProductNode_Float419: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float419weight,vb2,ProductNode_Float419Output_532);

SumNode_Float113: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float133Output_164,ProductNode_Float132Output_163,SumNode_Float113Output_533);

ProductNode_Float420: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float31Output_165,ProductNode_Float131Output_162,ProductNode_Float420Output_534);

SumNode_Float114: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float134Output_166,ProductNode_Float127Output_157,SumNode_Float114Output_535);

ProductNode_Float421: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb13,SumNode_Float32Output_167,ProductNode_Float421Output_536);

ProductNode_Float422: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float422weight,ProductNode_Float135Output_168,ProductNode_Float422Output_537);

SumNode_Float115: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float136Output_169,ProductNode_Float120Output_148,SumNode_Float115Output_538);

ProductNode_Float423: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v10,SumNode_Float33Output_170,ProductNode_Float423Output_539);

ProductNode_Float424: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float424weight,v1,ProductNode_Float424Output_540);

ProductNode_Float425: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float425weight,vb1,ProductNode_Float425Output_541);

SumNode_Float116: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float139Output_173,ProductNode_Float138Output_172,SumNode_Float116Output_542);

ProductNode_Float426: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v9,SumNode_Float34Output_174,ProductNode_Float426Output_543);

ProductNode_Float427: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float427weight,ProductNode_Float140Output_175,ProductNode_Float427Output_544);

ProductNode_Float428: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float428weight,ProductNode_Float141Output_176,ProductNode_Float428Output_545);

ProductNode_Float429: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float429weight,v1,ProductNode_Float429Output_546);

ProductNode_Float430: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float430weight,vb1,ProductNode_Float430Output_547);

SumNode_Float117: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float144Output_179,ProductNode_Float143Output_178,SumNode_Float117Output_548);

ProductNode_Float431: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb9,SumNode_Float35Output_180,ProductNode_Float431Output_549);

ProductNode_Float432: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float432weight,ProductNode_Float145Output_181,ProductNode_Float432Output_550);

ProductNode_Float433: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float433weight,ProductNode_Float146Output_182,ProductNode_Float433Output_551);

SumNode_Float118: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float147Output_183,ProductNode_Float142Output_177,SumNode_Float118Output_552);

ProductNode_Float434: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float36Output_184,ProductNode_Float137Output_171,ProductNode_Float434Output_553);

ProductNode_Float435: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float435weight,v11,ProductNode_Float435Output_554);

ProductNode_Float436: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float436weight,vb11,ProductNode_Float436Output_555);

SumNode_Float119: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float106Output_129,ProductNode_Float105Output_128,SumNode_Float119Output_556);

ProductNode_Float437: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v12,SumNode_Float23Output_130,ProductNode_Float437Output_557);

ProductNode_Float438: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float438weight,ProductNode_Float107Output_131,ProductNode_Float438Output_558);

ProductNode_Float439: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float439weight,v2,ProductNode_Float439Output_559);

ProductNode_Float440: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float440weight,vb2,ProductNode_Float440Output_560);

SumNode_Float120: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float110Output_134,ProductNode_Float109Output_133,SumNode_Float120Output_561);

ProductNode_Float441: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float24Output_135,ProductNode_Float108Output_132,ProductNode_Float441Output_562);

ProductNode_Float442: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float442weight,v11,ProductNode_Float442Output_563);

ProductNode_Float443: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float443weight,vb11,ProductNode_Float443Output_564);

SumNode_Float121: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float113Output_138,ProductNode_Float112Output_137,SumNode_Float121Output_565);

ProductNode_Float444: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb12,SumNode_Float25Output_139,ProductNode_Float444Output_566);

ProductNode_Float445: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float445weight,ProductNode_Float114Output_140,ProductNode_Float445Output_567);

ProductNode_Float446: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float446weight,v2,ProductNode_Float446Output_568);

ProductNode_Float447: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float447weight,vb2,ProductNode_Float447Output_569);

SumNode_Float122: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float117Output_143,ProductNode_Float116Output_142,SumNode_Float122Output_570);

ProductNode_Float448: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float26Output_144,ProductNode_Float115Output_141,ProductNode_Float448Output_571);

SumNode_Float123: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float118Output_145,ProductNode_Float111Output_136,SumNode_Float123Output_572);

ProductNode_Float449: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v13,SumNode_Float27Output_146,ProductNode_Float449Output_573);

ProductNode_Float450: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float450weight,ProductNode_Float119Output_147,ProductNode_Float450Output_574);

ProductNode_Float451: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float451weight,v11,ProductNode_Float451Output_575);

ProductNode_Float452: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float452weight,vb11,ProductNode_Float452Output_576);

SumNode_Float124: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float122Output_150,ProductNode_Float121Output_149,SumNode_Float124Output_577);

ProductNode_Float453: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v12,SumNode_Float28Output_151,ProductNode_Float453Output_578);

ProductNode_Float454: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float454weight,ProductNode_Float123Output_152,ProductNode_Float454Output_579);

ProductNode_Float455: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float455weight,v2,ProductNode_Float455Output_580);

ProductNode_Float456: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float456weight,vb2,ProductNode_Float456Output_581);

SumNode_Float125: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float126Output_155,ProductNode_Float125Output_154,SumNode_Float125Output_582);

ProductNode_Float457: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float29Output_156,ProductNode_Float124Output_153,ProductNode_Float457Output_583);

ProductNode_Float458: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float458weight,v11,ProductNode_Float458Output_584);

ProductNode_Float459: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float459weight,vb11,ProductNode_Float459Output_585);

SumNode_Float126: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float129Output_159,ProductNode_Float128Output_158,SumNode_Float126Output_586);

ProductNode_Float460: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb12,SumNode_Float30Output_160,ProductNode_Float460Output_587);

ProductNode_Float461: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float461weight,ProductNode_Float130Output_161,ProductNode_Float461Output_588);

ProductNode_Float462: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float462weight,v2,ProductNode_Float462Output_589);

ProductNode_Float463: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float463weight,vb2,ProductNode_Float463Output_590);

SumNode_Float127: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float133Output_164,ProductNode_Float132Output_163,SumNode_Float127Output_591);

ProductNode_Float464: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float31Output_165,ProductNode_Float131Output_162,ProductNode_Float464Output_592);

SumNode_Float128: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float134Output_166,ProductNode_Float127Output_157,SumNode_Float128Output_593);

ProductNode_Float465: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb13,SumNode_Float32Output_167,ProductNode_Float465Output_594);

ProductNode_Float466: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float466weight,ProductNode_Float135Output_168,ProductNode_Float466Output_595);

SumNode_Float129: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float180Output_227,ProductNode_Float164Output_206,SumNode_Float129Output_596);

ProductNode_Float467: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb10,SumNode_Float47Output_228,ProductNode_Float467Output_597);

ProductNode_Float468: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float468weight,v1,ProductNode_Float468Output_598);

ProductNode_Float469: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float469weight,vb1,ProductNode_Float469Output_599);

SumNode_Float130: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float183Output_231,ProductNode_Float182Output_230,SumNode_Float130Output_600);

ProductNode_Float470: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v9,SumNode_Float48Output_232,ProductNode_Float470Output_601);

ProductNode_Float471: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float471weight,ProductNode_Float184Output_233,ProductNode_Float471Output_602);

ProductNode_Float472: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float472weight,ProductNode_Float185Output_234,ProductNode_Float472Output_603);

ProductNode_Float473: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float473weight,v1,ProductNode_Float473Output_604);

ProductNode_Float474: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float474weight,vb1,ProductNode_Float474Output_605);

SumNode_Float131: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float188Output_237,ProductNode_Float187Output_236,SumNode_Float131Output_606);

ProductNode_Float475: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb9,SumNode_Float49Output_238,ProductNode_Float475Output_607);

ProductNode_Float476: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float476weight,ProductNode_Float189Output_239,ProductNode_Float476Output_608);

ProductNode_Float477: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float477weight,ProductNode_Float190Output_240,ProductNode_Float477Output_609);

SumNode_Float132: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float191Output_241,ProductNode_Float186Output_235,SumNode_Float132Output_610);

ProductNode_Float478: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float50Output_242,ProductNode_Float181Output_229,ProductNode_Float478Output_611);

SumNode_Float133: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float192Output_243,ProductNode_Float148Output_185,SumNode_Float133Output_612);

ProductNode_Float479: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v15,SumNode_Float51Output_244,ProductNode_Float479Output_613);

ProductNode_Float480: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float480weight,ProductNode_Float193Output_245,ProductNode_Float480Output_614);

ProductNode_Float481: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float481weight,v11,ProductNode_Float481Output_615);

ProductNode_Float482: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float482weight,vb11,ProductNode_Float482Output_616);

SumNode_Float134: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float106Output_129,ProductNode_Float105Output_128,SumNode_Float134Output_617);

ProductNode_Float483: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v12,SumNode_Float23Output_130,ProductNode_Float483Output_618);

ProductNode_Float484: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float484weight,ProductNode_Float107Output_131,ProductNode_Float484Output_619);

ProductNode_Float485: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float485weight,v2,ProductNode_Float485Output_620);

ProductNode_Float486: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float486weight,vb2,ProductNode_Float486Output_621);

SumNode_Float135: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float200Output_253,ProductNode_Float199Output_252,SumNode_Float135Output_622);

ProductNode_Float487: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float53Output_254,ProductNode_Float108Output_132,ProductNode_Float487Output_623);

ProductNode_Float488: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float488weight,v11,ProductNode_Float488Output_624);

ProductNode_Float489: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float489weight,vb11,ProductNode_Float489Output_625);

SumNode_Float136: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float113Output_138,ProductNode_Float112Output_137,SumNode_Float136Output_626);

ProductNode_Float490: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb12,SumNode_Float25Output_139,ProductNode_Float490Output_627);

ProductNode_Float491: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float491weight,ProductNode_Float114Output_140,ProductNode_Float491Output_628);

ProductNode_Float492: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float492weight,v2,ProductNode_Float492Output_629);

ProductNode_Float493: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float493weight,vb2,ProductNode_Float493Output_630);

SumNode_Float137: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float207Output_262,ProductNode_Float206Output_261,SumNode_Float137Output_631);

ProductNode_Float494: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float55Output_263,ProductNode_Float115Output_141,ProductNode_Float494Output_632);

SumNode_Float138: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float208Output_264,ProductNode_Float201Output_255,SumNode_Float138Output_633);

ProductNode_Float495: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v13,SumNode_Float56Output_265,ProductNode_Float495Output_634);

ProductNode_Float496: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float496weight,ProductNode_Float209Output_266,ProductNode_Float496Output_635);

ProductNode_Float497: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float497weight,v11,ProductNode_Float497Output_636);

ProductNode_Float498: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float498weight,vb11,ProductNode_Float498Output_637);

SumNode_Float139: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float122Output_150,ProductNode_Float121Output_149,SumNode_Float139Output_638);

ProductNode_Float499: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v12,SumNode_Float28Output_151,ProductNode_Float499Output_639);

ProductNode_Float500: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float500weight,ProductNode_Float123Output_152,ProductNode_Float500Output_640);

ProductNode_Float501: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float501weight,v2,ProductNode_Float501Output_641);

ProductNode_Float502: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float502weight,vb2,ProductNode_Float502Output_642);

SumNode_Float140: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float216Output_274,ProductNode_Float215Output_273,SumNode_Float140Output_643);

ProductNode_Float503: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float58Output_275,ProductNode_Float124Output_153,ProductNode_Float503Output_644);

ProductNode_Float504: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float504weight,v11,ProductNode_Float504Output_645);

ProductNode_Float505: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float505weight,vb11,ProductNode_Float505Output_646);

SumNode_Float141: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float129Output_159,ProductNode_Float128Output_158,SumNode_Float141Output_647);

ProductNode_Float506: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb12,SumNode_Float30Output_160,ProductNode_Float506Output_648);

ProductNode_Float507: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float507weight,ProductNode_Float130Output_161,ProductNode_Float507Output_649);

ProductNode_Float508: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float508weight,v2,ProductNode_Float508Output_650);

ProductNode_Float509: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float509weight,vb2,ProductNode_Float509Output_651);

SumNode_Float142: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float223Output_283,ProductNode_Float222Output_282,SumNode_Float142Output_652);

ProductNode_Float510: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float60Output_284,ProductNode_Float131Output_162,ProductNode_Float510Output_653);

SumNode_Float143: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float224Output_285,ProductNode_Float217Output_276,SumNode_Float143Output_654);

ProductNode_Float511: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb13,SumNode_Float61Output_286,ProductNode_Float511Output_655);

ProductNode_Float512: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float512weight,ProductNode_Float225Output_287,ProductNode_Float512Output_656);

SumNode_Float144: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float226Output_288,ProductNode_Float210Output_267,SumNode_Float144Output_657);

ProductNode_Float513: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v10,SumNode_Float62Output_289,ProductNode_Float513Output_658);

ProductNode_Float514: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float514weight,v1,ProductNode_Float514Output_659);

ProductNode_Float515: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float515weight,vb1,ProductNode_Float515Output_660);

SumNode_Float145: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float139Output_173,ProductNode_Float138Output_172,SumNode_Float145Output_661);

ProductNode_Float516: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v9,SumNode_Float34Output_174,ProductNode_Float516Output_662);

ProductNode_Float517: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float517weight,ProductNode_Float140Output_175,ProductNode_Float517Output_663);

ProductNode_Float518: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float518weight,ProductNode_Float231Output_295,ProductNode_Float518Output_664);

ProductNode_Float519: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float519weight,v1,ProductNode_Float519Output_665);

ProductNode_Float520: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float520weight,vb1,ProductNode_Float520Output_666);

SumNode_Float146: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float144Output_179,ProductNode_Float143Output_178,SumNode_Float146Output_667);

ProductNode_Float521: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb9,SumNode_Float35Output_180,ProductNode_Float521Output_668);

ProductNode_Float522: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float522weight,ProductNode_Float145Output_181,ProductNode_Float522Output_669);

ProductNode_Float523: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float523weight,ProductNode_Float236Output_301,ProductNode_Float523Output_670);

SumNode_Float147: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float237Output_302,ProductNode_Float232Output_296,SumNode_Float147Output_671);

ProductNode_Float524: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float65Output_303,ProductNode_Float227Output_290,ProductNode_Float524Output_672);

ProductNode_Float525: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float525weight,v11,ProductNode_Float525Output_673);

ProductNode_Float526: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float526weight,vb11,ProductNode_Float526Output_674);

SumNode_Float148: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float106Output_129,ProductNode_Float105Output_128,SumNode_Float148Output_675);

ProductNode_Float527: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v12,SumNode_Float23Output_130,ProductNode_Float527Output_676);

ProductNode_Float528: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float528weight,ProductNode_Float107Output_131,ProductNode_Float528Output_677);

ProductNode_Float529: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float529weight,v2,ProductNode_Float529Output_678);

ProductNode_Float530: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float530weight,vb2,ProductNode_Float530Output_679);

SumNode_Float149: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float200Output_253,ProductNode_Float199Output_252,SumNode_Float149Output_680);

ProductNode_Float531: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float53Output_254,ProductNode_Float108Output_132,ProductNode_Float531Output_681);

ProductNode_Float532: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float532weight,v11,ProductNode_Float532Output_682);

ProductNode_Float533: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float533weight,vb11,ProductNode_Float533Output_683);

SumNode_Float150: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float113Output_138,ProductNode_Float112Output_137,SumNode_Float150Output_684);

ProductNode_Float534: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb12,SumNode_Float25Output_139,ProductNode_Float534Output_685);

ProductNode_Float535: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float535weight,ProductNode_Float114Output_140,ProductNode_Float535Output_686);

ProductNode_Float536: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float536weight,v2,ProductNode_Float536Output_687);

ProductNode_Float537: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float537weight,vb2,ProductNode_Float537Output_688);

SumNode_Float151: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float207Output_262,ProductNode_Float206Output_261,SumNode_Float151Output_689);

ProductNode_Float538: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float55Output_263,ProductNode_Float115Output_141,ProductNode_Float538Output_690);

SumNode_Float152: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float208Output_264,ProductNode_Float201Output_255,SumNode_Float152Output_691);

ProductNode_Float539: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v13,SumNode_Float56Output_265,ProductNode_Float539Output_692);

ProductNode_Float540: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float540weight,ProductNode_Float209Output_266,ProductNode_Float540Output_693);

ProductNode_Float541: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float541weight,v11,ProductNode_Float541Output_694);

ProductNode_Float542: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float542weight,vb11,ProductNode_Float542Output_695);

SumNode_Float153: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float122Output_150,ProductNode_Float121Output_149,SumNode_Float153Output_696);

ProductNode_Float543: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v12,SumNode_Float28Output_151,ProductNode_Float543Output_697);

ProductNode_Float544: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float544weight,ProductNode_Float123Output_152,ProductNode_Float544Output_698);

ProductNode_Float545: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float545weight,v2,ProductNode_Float545Output_699);

ProductNode_Float546: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float546weight,vb2,ProductNode_Float546Output_700);

SumNode_Float154: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float216Output_274,ProductNode_Float215Output_273,SumNode_Float154Output_701);

ProductNode_Float547: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float58Output_275,ProductNode_Float124Output_153,ProductNode_Float547Output_702);

ProductNode_Float548: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float548weight,v11,ProductNode_Float548Output_703);

ProductNode_Float549: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float549weight,vb11,ProductNode_Float549Output_704);

SumNode_Float155: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float129Output_159,ProductNode_Float128Output_158,SumNode_Float155Output_705);

ProductNode_Float550: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb12,SumNode_Float30Output_160,ProductNode_Float550Output_706);

ProductNode_Float551: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float551weight,ProductNode_Float130Output_161,ProductNode_Float551Output_707);

ProductNode_Float552: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float552weight,v2,ProductNode_Float552Output_708);

ProductNode_Float553: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float553weight,vb2,ProductNode_Float553Output_709);

SumNode_Float156: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float223Output_283,ProductNode_Float222Output_282,SumNode_Float156Output_710);

ProductNode_Float554: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float60Output_284,ProductNode_Float131Output_162,ProductNode_Float554Output_711);

SumNode_Float157: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float224Output_285,ProductNode_Float217Output_276,SumNode_Float157Output_712);

ProductNode_Float555: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb13,SumNode_Float61Output_286,ProductNode_Float555Output_713);

ProductNode_Float556: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float556weight,ProductNode_Float225Output_287,ProductNode_Float556Output_714);

SumNode_Float158: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float270Output_346,ProductNode_Float254Output_325,SumNode_Float158Output_715);

ProductNode_Float557: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb10,SumNode_Float76Output_347,ProductNode_Float557Output_716);

ProductNode_Float558: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float558weight,v1,ProductNode_Float558Output_717);

ProductNode_Float559: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float559weight,vb1,ProductNode_Float559Output_718);

SumNode_Float159: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float183Output_231,ProductNode_Float182Output_230,SumNode_Float159Output_719);

ProductNode_Float560: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v9,SumNode_Float48Output_232,ProductNode_Float560Output_720);

ProductNode_Float561: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float561weight,ProductNode_Float184Output_233,ProductNode_Float561Output_721);

ProductNode_Float562: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float562weight,ProductNode_Float275Output_353,ProductNode_Float562Output_722);

ProductNode_Float563: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float563weight,v1,ProductNode_Float563Output_723);

ProductNode_Float564: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float564weight,vb1,ProductNode_Float564Output_724);

SumNode_Float160: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float188Output_237,ProductNode_Float187Output_236,SumNode_Float160Output_725);

ProductNode_Float565: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb9,SumNode_Float49Output_238,ProductNode_Float565Output_726);

ProductNode_Float566: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float566weight,ProductNode_Float189Output_239,ProductNode_Float566Output_727);

ProductNode_Float567: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float567weight,ProductNode_Float280Output_359,ProductNode_Float567Output_728);

SumNode_Float161: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float281Output_360,ProductNode_Float276Output_354,SumNode_Float161Output_729);

ProductNode_Float568: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float79Output_361,ProductNode_Float271Output_348,ProductNode_Float568Output_730);

SumNode_Float162: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float282Output_362,ProductNode_Float238Output_304,SumNode_Float162Output_731);

ProductNode_Float569: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb15,SumNode_Float80Output_363,ProductNode_Float569Output_732);

ProductNode_Float570: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float570weight,ProductNode_Float283Output_364,ProductNode_Float570Output_733);

SumNode_Float163: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float570Output_733,ProductNode_Float480Output_614,SumNode_Float163Output_734);

ProductNode_Float571: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float163Output_734,ProductNode_Float390Output_495,ProductNode_Float571Output_735);

SumNode_Float164: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float571Output_735,ProductNode_Float285Output_367,SumNode_Float164Output_736);

ProductNode_Float572: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v6,SumNode_Float164Output_736,ProductNode_Float572Output_737);

ProductNode_Float573: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float573weight,v4,ProductNode_Float573Output_738);

ProductNode_Float574: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float574weight,v8,ProductNode_Float574Output_739);

ProductNode_Float575: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float575weight,vb8,ProductNode_Float575Output_740);

SumNode_Float165: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2Output_2,ProductNode_Float1Output_1,SumNode_Float165Output_741);

ProductNode_Float576: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v7,SumNode_Float0Output_3,ProductNode_Float576Output_742);

ProductNode_Float577: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float577weight,v3,ProductNode_Float577Output_743);

ProductNode_Float578: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float578weight,ProductNode_Float4Output_5,ProductNode_Float578Output_744);

ProductNode_Float579: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float579weight,ProductNode_Float5Output_6,ProductNode_Float579Output_745);

ProductNode_Float580: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float580weight,vb3,ProductNode_Float580Output_746);

ProductNode_Float581: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float581weight,ProductNode_Float7Output_8,ProductNode_Float581Output_747);

ProductNode_Float582: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float582weight,ProductNode_Float8Output_9,ProductNode_Float582Output_748);

SumNode_Float166: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float9Output_10,ProductNode_Float6Output_7,SumNode_Float166Output_749);

ProductNode_Float583: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float1Output_11,ProductNode_Float3Output_4,ProductNode_Float583Output_750);

ProductNode_Float584: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float584weight,ProductNode_Float10Output_12,ProductNode_Float584Output_751);

ProductNode_Float585: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float585weight,v8,ProductNode_Float585Output_752);

ProductNode_Float586: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float586weight,vb8,ProductNode_Float586Output_753);

SumNode_Float167: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float13Output_15,ProductNode_Float12Output_14,SumNode_Float167Output_754);

ProductNode_Float587: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb7,SumNode_Float2Output_16,ProductNode_Float587Output_755);

ProductNode_Float588: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float588weight,v3,ProductNode_Float588Output_756);

ProductNode_Float589: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float589weight,ProductNode_Float4Output_5,ProductNode_Float589Output_757);

ProductNode_Float590: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float590weight,ProductNode_Float16Output_19,ProductNode_Float590Output_758);

ProductNode_Float591: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float591weight,vb3,ProductNode_Float591Output_759);

ProductNode_Float592: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float592weight,ProductNode_Float7Output_8,ProductNode_Float592Output_760);

ProductNode_Float593: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float593weight,ProductNode_Float19Output_22,ProductNode_Float593Output_761);

SumNode_Float168: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float20Output_23,ProductNode_Float17Output_20,SumNode_Float168Output_762);

ProductNode_Float594: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float3Output_24,ProductNode_Float14Output_17,ProductNode_Float594Output_763);

ProductNode_Float595: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float595weight,ProductNode_Float21Output_25,ProductNode_Float595Output_764);

SumNode_Float169: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float595Output_764,ProductNode_Float584Output_751,SumNode_Float169Output_765);

ProductNode_Float596: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float169Output_765,ProductNode_Float0Output_0,ProductNode_Float596Output_766);

ProductNode_Float597: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float597weight,ProductNode_Float596Output_766,ProductNode_Float597Output_767);

ProductNode_Float598: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float598weight,vb4,ProductNode_Float598Output_768);

ProductNode_Float599: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float599weight,v8,ProductNode_Float599Output_769);

ProductNode_Float600: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float600weight,vb8,ProductNode_Float600Output_770);

SumNode_Float170: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float27Output_32,ProductNode_Float26Output_31,SumNode_Float170Output_771);

ProductNode_Float601: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v7,SumNode_Float5Output_33,ProductNode_Float601Output_772);

ProductNode_Float602: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float602weight,v3,ProductNode_Float602Output_773);

ProductNode_Float603: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float603weight,ProductNode_Float29Output_35,ProductNode_Float603Output_774);

ProductNode_Float604: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float604weight,ProductNode_Float30Output_36,ProductNode_Float604Output_775);

ProductNode_Float605: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float605weight,vb3,ProductNode_Float605Output_776);

ProductNode_Float606: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float606weight,ProductNode_Float32Output_38,ProductNode_Float606Output_777);

ProductNode_Float607: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float607weight,ProductNode_Float33Output_39,ProductNode_Float607Output_778);

SumNode_Float171: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float34Output_40,ProductNode_Float31Output_37,SumNode_Float171Output_779);

ProductNode_Float608: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float6Output_41,ProductNode_Float28Output_34,ProductNode_Float608Output_780);

ProductNode_Float609: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float609weight,ProductNode_Float35Output_42,ProductNode_Float609Output_781);

ProductNode_Float610: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float610weight,v8,ProductNode_Float610Output_782);

ProductNode_Float611: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float611weight,vb8,ProductNode_Float611Output_783);

SumNode_Float172: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float38Output_45,ProductNode_Float37Output_44,SumNode_Float172Output_784);

ProductNode_Float612: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb7,SumNode_Float7Output_46,ProductNode_Float612Output_785);

ProductNode_Float613: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float613weight,v3,ProductNode_Float613Output_786);

ProductNode_Float614: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float614weight,ProductNode_Float29Output_35,ProductNode_Float614Output_787);

ProductNode_Float615: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float615weight,ProductNode_Float41Output_49,ProductNode_Float615Output_788);

ProductNode_Float616: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float616weight,vb3,ProductNode_Float616Output_789);

ProductNode_Float617: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float617weight,ProductNode_Float32Output_38,ProductNode_Float617Output_790);

ProductNode_Float618: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float618weight,ProductNode_Float44Output_52,ProductNode_Float618Output_791);

SumNode_Float173: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float45Output_53,ProductNode_Float42Output_50,SumNode_Float173Output_792);

ProductNode_Float619: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float8Output_54,ProductNode_Float39Output_47,ProductNode_Float619Output_793);

ProductNode_Float620: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float620weight,ProductNode_Float46Output_55,ProductNode_Float620Output_794);

SumNode_Float174: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float620Output_794,ProductNode_Float609Output_781,SumNode_Float174Output_795);

ProductNode_Float621: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float174Output_795,ProductNode_Float25Output_30,ProductNode_Float621Output_796);

ProductNode_Float622: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float622weight,ProductNode_Float621Output_796,ProductNode_Float622Output_797);

SumNode_Float175: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float622Output_797,ProductNode_Float597Output_767,SumNode_Float175Output_798);

ProductNode_Float623: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v5,SumNode_Float175Output_798,ProductNode_Float623Output_799);

ProductNode_Float624: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float624weight,ProductNode_Float623Output_799,ProductNode_Float624Output_800);

ProductNode_Float625: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float625weight,v4,ProductNode_Float625Output_801);

ProductNode_Float626: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float626weight,v8,ProductNode_Float626Output_802);

ProductNode_Float627: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float627weight,vb8,ProductNode_Float627Output_803);

SumNode_Float176: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float54Output_65,ProductNode_Float53Output_64,SumNode_Float176Output_804);

ProductNode_Float628: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v7,SumNode_Float11Output_66,ProductNode_Float628Output_805);

ProductNode_Float629: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float629weight,v3,ProductNode_Float629Output_806);

ProductNode_Float630: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float630weight,ProductNode_Float4Output_5,ProductNode_Float630Output_807);

ProductNode_Float631: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float631weight,ProductNode_Float5Output_6,ProductNode_Float631Output_808);

ProductNode_Float632: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float632weight,vb3,ProductNode_Float632Output_809);

ProductNode_Float633: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float633weight,ProductNode_Float7Output_8,ProductNode_Float633Output_810);

ProductNode_Float634: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float634weight,ProductNode_Float8Output_9,ProductNode_Float634Output_811);

SumNode_Float177: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float61Output_73,ProductNode_Float58Output_70,SumNode_Float177Output_812);

ProductNode_Float635: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float12Output_74,ProductNode_Float55Output_67,ProductNode_Float635Output_813);

ProductNode_Float636: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float636weight,ProductNode_Float62Output_75,ProductNode_Float636Output_814);

ProductNode_Float637: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float637weight,v8,ProductNode_Float637Output_815);

ProductNode_Float638: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float638weight,vb8,ProductNode_Float638Output_816);

SumNode_Float178: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float65Output_78,ProductNode_Float64Output_77,SumNode_Float178Output_817);

ProductNode_Float639: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb7,SumNode_Float13Output_79,ProductNode_Float639Output_818);

ProductNode_Float640: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float640weight,v3,ProductNode_Float640Output_819);

ProductNode_Float641: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float641weight,ProductNode_Float4Output_5,ProductNode_Float641Output_820);

ProductNode_Float642: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float642weight,ProductNode_Float16Output_19,ProductNode_Float642Output_821);

ProductNode_Float643: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float643weight,vb3,ProductNode_Float643Output_822);

ProductNode_Float644: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float644weight,ProductNode_Float7Output_8,ProductNode_Float644Output_823);

ProductNode_Float645: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float645weight,ProductNode_Float19Output_22,ProductNode_Float645Output_824);

SumNode_Float179: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float72Output_86,ProductNode_Float69Output_83,SumNode_Float179Output_825);

ProductNode_Float646: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float14Output_87,ProductNode_Float66Output_80,ProductNode_Float646Output_826);

ProductNode_Float647: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float647weight,ProductNode_Float73Output_88,ProductNode_Float647Output_827);

SumNode_Float180: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float647Output_827,ProductNode_Float636Output_814,SumNode_Float180Output_828);

ProductNode_Float648: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float180Output_828,ProductNode_Float0Output_0,ProductNode_Float648Output_829);

ProductNode_Float649: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float649weight,ProductNode_Float648Output_829,ProductNode_Float649Output_830);

ProductNode_Float650: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float650weight,vb4,ProductNode_Float650Output_831);

ProductNode_Float651: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float651weight,v8,ProductNode_Float651Output_832);

ProductNode_Float652: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float652weight,vb8,ProductNode_Float652Output_833);

SumNode_Float181: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float79Output_95,ProductNode_Float78Output_94,SumNode_Float181Output_834);

ProductNode_Float653: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v7,SumNode_Float16Output_96,ProductNode_Float653Output_835);

ProductNode_Float654: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float654weight,v3,ProductNode_Float654Output_836);

ProductNode_Float655: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float655weight,ProductNode_Float29Output_35,ProductNode_Float655Output_837);

ProductNode_Float656: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float656weight,ProductNode_Float30Output_36,ProductNode_Float656Output_838);

ProductNode_Float657: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float657weight,vb3,ProductNode_Float657Output_839);

ProductNode_Float658: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float658weight,ProductNode_Float32Output_38,ProductNode_Float658Output_840);

ProductNode_Float659: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float659weight,ProductNode_Float33Output_39,ProductNode_Float659Output_841);

SumNode_Float182: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float86Output_103,ProductNode_Float83Output_100,SumNode_Float182Output_842);

ProductNode_Float660: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float17Output_104,ProductNode_Float80Output_97,ProductNode_Float660Output_843);

ProductNode_Float661: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float661weight,ProductNode_Float87Output_105,ProductNode_Float661Output_844);

ProductNode_Float662: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float662weight,v8,ProductNode_Float662Output_845);

ProductNode_Float663: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float663weight,vb8,ProductNode_Float663Output_846);

SumNode_Float183: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float90Output_108,ProductNode_Float89Output_107,SumNode_Float183Output_847);

ProductNode_Float664: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb7,SumNode_Float18Output_109,ProductNode_Float664Output_848);

ProductNode_Float665: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float665weight,v3,ProductNode_Float665Output_849);

ProductNode_Float666: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float666weight,ProductNode_Float29Output_35,ProductNode_Float666Output_850);

ProductNode_Float667: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float667weight,ProductNode_Float41Output_49,ProductNode_Float667Output_851);

ProductNode_Float668: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float668weight,vb3,ProductNode_Float668Output_852);

ProductNode_Float669: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float669weight,ProductNode_Float32Output_38,ProductNode_Float669Output_853);

ProductNode_Float670: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float670weight,ProductNode_Float44Output_52,ProductNode_Float670Output_854);

SumNode_Float184: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float97Output_116,ProductNode_Float94Output_113,SumNode_Float184Output_855);

ProductNode_Float671: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float19Output_117,ProductNode_Float91Output_110,ProductNode_Float671Output_856);

ProductNode_Float672: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float672weight,ProductNode_Float98Output_118,ProductNode_Float672Output_857);

SumNode_Float185: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float672Output_857,ProductNode_Float661Output_844,SumNode_Float185Output_858);

ProductNode_Float673: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float185Output_858,ProductNode_Float25Output_30,ProductNode_Float673Output_859);

ProductNode_Float674: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float674weight,ProductNode_Float673Output_859,ProductNode_Float674Output_860);

SumNode_Float186: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float674Output_860,ProductNode_Float649Output_830,SumNode_Float186Output_861);

ProductNode_Float675: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb5,SumNode_Float186Output_861,ProductNode_Float675Output_862);

ProductNode_Float676: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float676weight,ProductNode_Float675Output_862,ProductNode_Float676Output_863);

SumNode_Float187: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float676Output_863,ProductNode_Float624Output_800,SumNode_Float187Output_864);

ProductNode_Float677: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v16,SumNode_Float187Output_864,ProductNode_Float677Output_865);

ProductNode_Float678: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float678weight,v11,ProductNode_Float678Output_866);

ProductNode_Float679: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float679weight,vb11,ProductNode_Float679Output_867);

SumNode_Float188: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float679Output_867,ProductNode_Float678Output_866,SumNode_Float188Output_868);

ProductNode_Float680: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v12,SumNode_Float188Output_868,ProductNode_Float680Output_869);

ProductNode_Float681: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float681weight,ProductNode_Float680Output_869,ProductNode_Float681Output_870);

ProductNode_Float682: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float682weight,v2,ProductNode_Float682Output_871);

ProductNode_Float683: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float683weight,vb2,ProductNode_Float683Output_872);

SumNode_Float189: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float110Output_134,ProductNode_Float109Output_133,SumNode_Float189Output_873);

ProductNode_Float684: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float24Output_135,ProductNode_Float681Output_870,ProductNode_Float684Output_874);

ProductNode_Float685: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float685weight,v11,ProductNode_Float685Output_875);

ProductNode_Float686: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float686weight,vb11,ProductNode_Float686Output_876);

SumNode_Float190: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float686Output_876,ProductNode_Float685Output_875,SumNode_Float190Output_877);

ProductNode_Float687: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb12,SumNode_Float190Output_877,ProductNode_Float687Output_878);

ProductNode_Float688: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float688weight,ProductNode_Float687Output_878,ProductNode_Float688Output_879);

ProductNode_Float689: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float689weight,v2,ProductNode_Float689Output_880);

ProductNode_Float690: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float690weight,vb2,ProductNode_Float690Output_881);

SumNode_Float191: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float117Output_143,ProductNode_Float116Output_142,SumNode_Float191Output_882);

ProductNode_Float691: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float26Output_144,ProductNode_Float688Output_879,ProductNode_Float691Output_883);

SumNode_Float192: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float691Output_883,ProductNode_Float684Output_874,SumNode_Float192Output_884);

ProductNode_Float692: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v13,SumNode_Float192Output_884,ProductNode_Float692Output_885);

ProductNode_Float693: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float693weight,ProductNode_Float692Output_885,ProductNode_Float693Output_886);

ProductNode_Float694: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float694weight,v11,ProductNode_Float694Output_887);

ProductNode_Float695: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float695weight,vb11,ProductNode_Float695Output_888);

SumNode_Float193: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float695Output_888,ProductNode_Float694Output_887,SumNode_Float193Output_889);

ProductNode_Float696: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v12,SumNode_Float193Output_889,ProductNode_Float696Output_890);

ProductNode_Float697: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float697weight,ProductNode_Float696Output_890,ProductNode_Float697Output_891);

ProductNode_Float698: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float698weight,v2,ProductNode_Float698Output_892);

ProductNode_Float699: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float699weight,vb2,ProductNode_Float699Output_893);

SumNode_Float194: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float126Output_155,ProductNode_Float125Output_154,SumNode_Float194Output_894);

ProductNode_Float700: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float29Output_156,ProductNode_Float697Output_891,ProductNode_Float700Output_895);

ProductNode_Float701: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float701weight,v11,ProductNode_Float701Output_896);

ProductNode_Float702: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float702weight,vb11,ProductNode_Float702Output_897);

SumNode_Float195: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float702Output_897,ProductNode_Float701Output_896,SumNode_Float195Output_898);

ProductNode_Float703: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb12,SumNode_Float195Output_898,ProductNode_Float703Output_899);

ProductNode_Float704: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float704weight,ProductNode_Float703Output_899,ProductNode_Float704Output_900);

ProductNode_Float705: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float705weight,v2,ProductNode_Float705Output_901);

ProductNode_Float706: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float706weight,vb2,ProductNode_Float706Output_902);

SumNode_Float196: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float133Output_164,ProductNode_Float132Output_163,SumNode_Float196Output_903);

ProductNode_Float707: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float31Output_165,ProductNode_Float704Output_900,ProductNode_Float707Output_904);

SumNode_Float197: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float707Output_904,ProductNode_Float700Output_895,SumNode_Float197Output_905);

ProductNode_Float708: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb13,SumNode_Float197Output_905,ProductNode_Float708Output_906);

ProductNode_Float709: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float709weight,ProductNode_Float708Output_906,ProductNode_Float709Output_907);

SumNode_Float198: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float709Output_907,ProductNode_Float693Output_886,SumNode_Float198Output_908);

ProductNode_Float710: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v10,SumNode_Float198Output_908,ProductNode_Float710Output_909);

ProductNode_Float711: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float711weight,v1,ProductNode_Float711Output_910);

ProductNode_Float712: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float712weight,vb1,ProductNode_Float712Output_911);

SumNode_Float199: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float139Output_173,ProductNode_Float138Output_172,SumNode_Float199Output_912);

ProductNode_Float713: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v9,SumNode_Float34Output_174,ProductNode_Float713Output_913);

ProductNode_Float714: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float714weight,ProductNode_Float140Output_175,ProductNode_Float714Output_914);

ProductNode_Float715: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float715weight,ProductNode_Float141Output_176,ProductNode_Float715Output_915);

ProductNode_Float716: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float716weight,v1,ProductNode_Float716Output_916);

ProductNode_Float717: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float717weight,vb1,ProductNode_Float717Output_917);

SumNode_Float200: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float144Output_179,ProductNode_Float143Output_178,SumNode_Float200Output_918);

ProductNode_Float718: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb9,SumNode_Float35Output_180,ProductNode_Float718Output_919);

ProductNode_Float719: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float719weight,ProductNode_Float145Output_181,ProductNode_Float719Output_920);

ProductNode_Float720: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float720weight,ProductNode_Float146Output_182,ProductNode_Float720Output_921);

SumNode_Float201: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float147Output_183,ProductNode_Float142Output_177,SumNode_Float201Output_922);

ProductNode_Float721: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float36Output_184,ProductNode_Float710Output_909,ProductNode_Float721Output_923);

ProductNode_Float722: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float722weight,v11,ProductNode_Float722Output_924);

ProductNode_Float723: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float723weight,vb11,ProductNode_Float723Output_925);

SumNode_Float202: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float679Output_867,ProductNode_Float678Output_866,SumNode_Float202Output_926);

ProductNode_Float724: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v12,SumNode_Float188Output_868,ProductNode_Float724Output_927);

ProductNode_Float725: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float725weight,ProductNode_Float680Output_869,ProductNode_Float725Output_928);

ProductNode_Float726: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float726weight,v2,ProductNode_Float726Output_929);

ProductNode_Float727: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float727weight,vb2,ProductNode_Float727Output_930);

SumNode_Float203: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float110Output_134,ProductNode_Float109Output_133,SumNode_Float203Output_931);

ProductNode_Float728: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float24Output_135,ProductNode_Float681Output_870,ProductNode_Float728Output_932);

ProductNode_Float729: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float729weight,v11,ProductNode_Float729Output_933);

ProductNode_Float730: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float730weight,vb11,ProductNode_Float730Output_934);

SumNode_Float204: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float686Output_876,ProductNode_Float685Output_875,SumNode_Float204Output_935);

ProductNode_Float731: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb12,SumNode_Float190Output_877,ProductNode_Float731Output_936);

ProductNode_Float732: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float732weight,ProductNode_Float687Output_878,ProductNode_Float732Output_937);

ProductNode_Float733: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float733weight,v2,ProductNode_Float733Output_938);

ProductNode_Float734: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float734weight,vb2,ProductNode_Float734Output_939);

SumNode_Float205: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float117Output_143,ProductNode_Float116Output_142,SumNode_Float205Output_940);

ProductNode_Float735: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float26Output_144,ProductNode_Float688Output_879,ProductNode_Float735Output_941);

SumNode_Float206: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float691Output_883,ProductNode_Float684Output_874,SumNode_Float206Output_942);

ProductNode_Float736: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v13,SumNode_Float192Output_884,ProductNode_Float736Output_943);

ProductNode_Float737: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float737weight,ProductNode_Float692Output_885,ProductNode_Float737Output_944);

ProductNode_Float738: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float738weight,v11,ProductNode_Float738Output_945);

ProductNode_Float739: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float739weight,vb11,ProductNode_Float739Output_946);

SumNode_Float207: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float695Output_888,ProductNode_Float694Output_887,SumNode_Float207Output_947);

ProductNode_Float740: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v12,SumNode_Float193Output_889,ProductNode_Float740Output_948);

ProductNode_Float741: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float741weight,ProductNode_Float696Output_890,ProductNode_Float741Output_949);

ProductNode_Float742: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float742weight,v2,ProductNode_Float742Output_950);

ProductNode_Float743: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float743weight,vb2,ProductNode_Float743Output_951);

SumNode_Float208: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float126Output_155,ProductNode_Float125Output_154,SumNode_Float208Output_952);

ProductNode_Float744: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float29Output_156,ProductNode_Float697Output_891,ProductNode_Float744Output_953);

ProductNode_Float745: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float745weight,v11,ProductNode_Float745Output_954);

ProductNode_Float746: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float746weight,vb11,ProductNode_Float746Output_955);

SumNode_Float209: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float702Output_897,ProductNode_Float701Output_896,SumNode_Float209Output_956);

ProductNode_Float747: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb12,SumNode_Float195Output_898,ProductNode_Float747Output_957);

ProductNode_Float748: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float748weight,ProductNode_Float703Output_899,ProductNode_Float748Output_958);

ProductNode_Float749: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float749weight,v2,ProductNode_Float749Output_959);

ProductNode_Float750: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float750weight,vb2,ProductNode_Float750Output_960);

SumNode_Float210: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float133Output_164,ProductNode_Float132Output_163,SumNode_Float210Output_961);

ProductNode_Float751: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float31Output_165,ProductNode_Float704Output_900,ProductNode_Float751Output_962);

SumNode_Float211: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float707Output_904,ProductNode_Float700Output_895,SumNode_Float211Output_963);

ProductNode_Float752: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb13,SumNode_Float197Output_905,ProductNode_Float752Output_964);

ProductNode_Float753: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float753weight,ProductNode_Float708Output_906,ProductNode_Float753Output_965);

SumNode_Float212: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float753Output_965,ProductNode_Float737Output_944,SumNode_Float212Output_966);

ProductNode_Float754: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb10,SumNode_Float212Output_966,ProductNode_Float754Output_967);

ProductNode_Float755: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float755weight,v1,ProductNode_Float755Output_968);

ProductNode_Float756: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float756weight,vb1,ProductNode_Float756Output_969);

SumNode_Float213: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float183Output_231,ProductNode_Float182Output_230,SumNode_Float213Output_970);

ProductNode_Float757: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v9,SumNode_Float48Output_232,ProductNode_Float757Output_971);

ProductNode_Float758: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float758weight,ProductNode_Float184Output_233,ProductNode_Float758Output_972);

ProductNode_Float759: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float759weight,ProductNode_Float185Output_234,ProductNode_Float759Output_973);

ProductNode_Float760: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float760weight,v1,ProductNode_Float760Output_974);

ProductNode_Float761: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float761weight,vb1,ProductNode_Float761Output_975);

SumNode_Float214: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float188Output_237,ProductNode_Float187Output_236,SumNode_Float214Output_976);

ProductNode_Float762: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb9,SumNode_Float49Output_238,ProductNode_Float762Output_977);

ProductNode_Float763: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float763weight,ProductNode_Float189Output_239,ProductNode_Float763Output_978);

ProductNode_Float764: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float764weight,ProductNode_Float190Output_240,ProductNode_Float764Output_979);

SumNode_Float215: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float191Output_241,ProductNode_Float186Output_235,SumNode_Float215Output_980);

ProductNode_Float765: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float50Output_242,ProductNode_Float754Output_967,ProductNode_Float765Output_981);

SumNode_Float216: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float765Output_981,ProductNode_Float721Output_923,SumNode_Float216Output_982);

ProductNode_Float766: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v15,SumNode_Float216Output_982,ProductNode_Float766Output_983);

ProductNode_Float767: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float767weight,ProductNode_Float766Output_983,ProductNode_Float767Output_984);

ProductNode_Float768: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float768weight,v11,ProductNode_Float768Output_985);

ProductNode_Float769: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float769weight,vb11,ProductNode_Float769Output_986);

SumNode_Float217: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float679Output_867,ProductNode_Float678Output_866,SumNode_Float217Output_987);

ProductNode_Float770: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v12,SumNode_Float188Output_868,ProductNode_Float770Output_988);

ProductNode_Float771: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float771weight,ProductNode_Float680Output_869,ProductNode_Float771Output_989);

ProductNode_Float772: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float772weight,v2,ProductNode_Float772Output_990);

ProductNode_Float773: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float773weight,vb2,ProductNode_Float773Output_991);

SumNode_Float218: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float200Output_253,ProductNode_Float199Output_252,SumNode_Float218Output_992);

ProductNode_Float774: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float53Output_254,ProductNode_Float681Output_870,ProductNode_Float774Output_993);

ProductNode_Float775: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float775weight,v11,ProductNode_Float775Output_994);

ProductNode_Float776: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float776weight,vb11,ProductNode_Float776Output_995);

SumNode_Float219: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float686Output_876,ProductNode_Float685Output_875,SumNode_Float219Output_996);

ProductNode_Float777: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb12,SumNode_Float190Output_877,ProductNode_Float777Output_997);

ProductNode_Float778: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float778weight,ProductNode_Float687Output_878,ProductNode_Float778Output_998);

ProductNode_Float779: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float779weight,v2,ProductNode_Float779Output_999);

ProductNode_Float780: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float780weight,vb2,ProductNode_Float780Output_1000);

SumNode_Float220: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float207Output_262,ProductNode_Float206Output_261,SumNode_Float220Output_1001);

ProductNode_Float781: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float55Output_263,ProductNode_Float688Output_879,ProductNode_Float781Output_1002);

SumNode_Float221: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float781Output_1002,ProductNode_Float774Output_993,SumNode_Float221Output_1003);

ProductNode_Float782: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v13,SumNode_Float221Output_1003,ProductNode_Float782Output_1004);

ProductNode_Float783: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float783weight,ProductNode_Float782Output_1004,ProductNode_Float783Output_1005);

ProductNode_Float784: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float784weight,v11,ProductNode_Float784Output_1006);

ProductNode_Float785: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float785weight,vb11,ProductNode_Float785Output_1007);

SumNode_Float222: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float695Output_888,ProductNode_Float694Output_887,SumNode_Float222Output_1008);

ProductNode_Float786: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v12,SumNode_Float193Output_889,ProductNode_Float786Output_1009);

ProductNode_Float787: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float787weight,ProductNode_Float696Output_890,ProductNode_Float787Output_1010);

ProductNode_Float788: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float788weight,v2,ProductNode_Float788Output_1011);

ProductNode_Float789: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float789weight,vb2,ProductNode_Float789Output_1012);

SumNode_Float223: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float216Output_274,ProductNode_Float215Output_273,SumNode_Float223Output_1013);

ProductNode_Float790: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float58Output_275,ProductNode_Float697Output_891,ProductNode_Float790Output_1014);

ProductNode_Float791: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float791weight,v11,ProductNode_Float791Output_1015);

ProductNode_Float792: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float792weight,vb11,ProductNode_Float792Output_1016);

SumNode_Float224: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float702Output_897,ProductNode_Float701Output_896,SumNode_Float224Output_1017);

ProductNode_Float793: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb12,SumNode_Float195Output_898,ProductNode_Float793Output_1018);

ProductNode_Float794: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float794weight,ProductNode_Float703Output_899,ProductNode_Float794Output_1019);

ProductNode_Float795: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float795weight,v2,ProductNode_Float795Output_1020);

ProductNode_Float796: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float796weight,vb2,ProductNode_Float796Output_1021);

SumNode_Float225: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float223Output_283,ProductNode_Float222Output_282,SumNode_Float225Output_1022);

ProductNode_Float797: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float60Output_284,ProductNode_Float704Output_900,ProductNode_Float797Output_1023);

SumNode_Float226: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float797Output_1023,ProductNode_Float790Output_1014,SumNode_Float226Output_1024);

ProductNode_Float798: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb13,SumNode_Float226Output_1024,ProductNode_Float798Output_1025);

ProductNode_Float799: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float799weight,ProductNode_Float798Output_1025,ProductNode_Float799Output_1026);

SumNode_Float227: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float799Output_1026,ProductNode_Float783Output_1005,SumNode_Float227Output_1027);

ProductNode_Float800: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v10,SumNode_Float227Output_1027,ProductNode_Float800Output_1028);

ProductNode_Float801: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float801weight,v1,ProductNode_Float801Output_1029);

ProductNode_Float802: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float802weight,vb1,ProductNode_Float802Output_1030);

SumNode_Float228: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float139Output_173,ProductNode_Float138Output_172,SumNode_Float228Output_1031);

ProductNode_Float803: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v9,SumNode_Float34Output_174,ProductNode_Float803Output_1032);

ProductNode_Float804: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float804weight,ProductNode_Float140Output_175,ProductNode_Float804Output_1033);

ProductNode_Float805: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float805weight,ProductNode_Float231Output_295,ProductNode_Float805Output_1034);

ProductNode_Float806: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float806weight,v1,ProductNode_Float806Output_1035);

ProductNode_Float807: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float807weight,vb1,ProductNode_Float807Output_1036);

SumNode_Float229: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float144Output_179,ProductNode_Float143Output_178,SumNode_Float229Output_1037);

ProductNode_Float808: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb9,SumNode_Float35Output_180,ProductNode_Float808Output_1038);

ProductNode_Float809: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float809weight,ProductNode_Float145Output_181,ProductNode_Float809Output_1039);

ProductNode_Float810: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float810weight,ProductNode_Float236Output_301,ProductNode_Float810Output_1040);

SumNode_Float230: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float237Output_302,ProductNode_Float232Output_296,SumNode_Float230Output_1041);

ProductNode_Float811: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float65Output_303,ProductNode_Float800Output_1028,ProductNode_Float811Output_1042);

ProductNode_Float812: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float812weight,v11,ProductNode_Float812Output_1043);

ProductNode_Float813: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float813weight,vb11,ProductNode_Float813Output_1044);

SumNode_Float231: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float679Output_867,ProductNode_Float678Output_866,SumNode_Float231Output_1045);

ProductNode_Float814: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v12,SumNode_Float188Output_868,ProductNode_Float814Output_1046);

ProductNode_Float815: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float815weight,ProductNode_Float680Output_869,ProductNode_Float815Output_1047);

ProductNode_Float816: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float816weight,v2,ProductNode_Float816Output_1048);

ProductNode_Float817: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float817weight,vb2,ProductNode_Float817Output_1049);

SumNode_Float232: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float200Output_253,ProductNode_Float199Output_252,SumNode_Float232Output_1050);

ProductNode_Float818: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float53Output_254,ProductNode_Float681Output_870,ProductNode_Float818Output_1051);

ProductNode_Float819: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float819weight,v11,ProductNode_Float819Output_1052);

ProductNode_Float820: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float820weight,vb11,ProductNode_Float820Output_1053);

SumNode_Float233: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float686Output_876,ProductNode_Float685Output_875,SumNode_Float233Output_1054);

ProductNode_Float821: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb12,SumNode_Float190Output_877,ProductNode_Float821Output_1055);

ProductNode_Float822: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float822weight,ProductNode_Float687Output_878,ProductNode_Float822Output_1056);

ProductNode_Float823: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float823weight,v2,ProductNode_Float823Output_1057);

ProductNode_Float824: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float824weight,vb2,ProductNode_Float824Output_1058);

SumNode_Float234: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float207Output_262,ProductNode_Float206Output_261,SumNode_Float234Output_1059);

ProductNode_Float825: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float55Output_263,ProductNode_Float688Output_879,ProductNode_Float825Output_1060);

SumNode_Float235: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float781Output_1002,ProductNode_Float774Output_993,SumNode_Float235Output_1061);

ProductNode_Float826: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v13,SumNode_Float221Output_1003,ProductNode_Float826Output_1062);

ProductNode_Float827: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float827weight,ProductNode_Float782Output_1004,ProductNode_Float827Output_1063);

ProductNode_Float828: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float828weight,v11,ProductNode_Float828Output_1064);

ProductNode_Float829: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float829weight,vb11,ProductNode_Float829Output_1065);

SumNode_Float236: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float695Output_888,ProductNode_Float694Output_887,SumNode_Float236Output_1066);

ProductNode_Float830: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v12,SumNode_Float193Output_889,ProductNode_Float830Output_1067);

ProductNode_Float831: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float831weight,ProductNode_Float696Output_890,ProductNode_Float831Output_1068);

ProductNode_Float832: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float832weight,v2,ProductNode_Float832Output_1069);

ProductNode_Float833: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float833weight,vb2,ProductNode_Float833Output_1070);

SumNode_Float237: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float216Output_274,ProductNode_Float215Output_273,SumNode_Float237Output_1071);

ProductNode_Float834: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float58Output_275,ProductNode_Float697Output_891,ProductNode_Float834Output_1072);

ProductNode_Float835: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float835weight,v11,ProductNode_Float835Output_1073);

ProductNode_Float836: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float836weight,vb11,ProductNode_Float836Output_1074);

SumNode_Float238: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float702Output_897,ProductNode_Float701Output_896,SumNode_Float238Output_1075);

ProductNode_Float837: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb12,SumNode_Float195Output_898,ProductNode_Float837Output_1076);

ProductNode_Float838: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float838weight,ProductNode_Float703Output_899,ProductNode_Float838Output_1077);

ProductNode_Float839: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float839weight,v2,ProductNode_Float839Output_1078);

ProductNode_Float840: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float840weight,vb2,ProductNode_Float840Output_1079);

SumNode_Float239: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float223Output_283,ProductNode_Float222Output_282,SumNode_Float239Output_1080);

ProductNode_Float841: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float60Output_284,ProductNode_Float704Output_900,ProductNode_Float841Output_1081);

SumNode_Float240: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float797Output_1023,ProductNode_Float790Output_1014,SumNode_Float240Output_1082);

ProductNode_Float842: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb13,SumNode_Float226Output_1024,ProductNode_Float842Output_1083);

ProductNode_Float843: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float843weight,ProductNode_Float798Output_1025,ProductNode_Float843Output_1084);

SumNode_Float241: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float843Output_1084,ProductNode_Float827Output_1063,SumNode_Float241Output_1085);

ProductNode_Float844: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb10,SumNode_Float241Output_1085,ProductNode_Float844Output_1086);

ProductNode_Float845: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float845weight,v1,ProductNode_Float845Output_1087);

ProductNode_Float846: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float846weight,vb1,ProductNode_Float846Output_1088);

SumNode_Float242: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float183Output_231,ProductNode_Float182Output_230,SumNode_Float242Output_1089);

ProductNode_Float847: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v9,SumNode_Float48Output_232,ProductNode_Float847Output_1090);

ProductNode_Float848: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float848weight,ProductNode_Float184Output_233,ProductNode_Float848Output_1091);

ProductNode_Float849: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float849weight,ProductNode_Float275Output_353,ProductNode_Float849Output_1092);

ProductNode_Float850: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float850weight,v1,ProductNode_Float850Output_1093);

ProductNode_Float851: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float851weight,vb1,ProductNode_Float851Output_1094);

SumNode_Float243: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float188Output_237,ProductNode_Float187Output_236,SumNode_Float243Output_1095);

ProductNode_Float852: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb9,SumNode_Float49Output_238,ProductNode_Float852Output_1096);

ProductNode_Float853: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float853weight,ProductNode_Float189Output_239,ProductNode_Float853Output_1097);

ProductNode_Float854: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float854weight,ProductNode_Float280Output_359,ProductNode_Float854Output_1098);

SumNode_Float244: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float281Output_360,ProductNode_Float276Output_354,SumNode_Float244Output_1099);

ProductNode_Float855: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float79Output_361,ProductNode_Float844Output_1086,ProductNode_Float855Output_1100);

SumNode_Float245: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float855Output_1100,ProductNode_Float811Output_1042,SumNode_Float245Output_1101);

ProductNode_Float856: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb15,SumNode_Float245Output_1101,ProductNode_Float856Output_1102);

ProductNode_Float857: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float857weight,ProductNode_Float856Output_1102,ProductNode_Float857Output_1103);

SumNode_Float246: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float857Output_1103,ProductNode_Float767Output_984,SumNode_Float246Output_1104);

ProductNode_Float858: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float246Output_1104,ProductNode_Float677Output_865,ProductNode_Float858Output_1105);

ProductNode_Float859: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float859weight,v4,ProductNode_Float859Output_1106);

ProductNode_Float860: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float860weight,v8,ProductNode_Float860Output_1107);

ProductNode_Float861: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float861weight,vb8,ProductNode_Float861Output_1108);

SumNode_Float247: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2Output_2,ProductNode_Float1Output_1,SumNode_Float247Output_1109);

ProductNode_Float862: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v7,SumNode_Float0Output_3,ProductNode_Float862Output_1110);

ProductNode_Float863: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float863weight,v3,ProductNode_Float863Output_1111);

ProductNode_Float864: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float864weight,ProductNode_Float4Output_5,ProductNode_Float864Output_1112);

ProductNode_Float865: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float865weight,ProductNode_Float5Output_6,ProductNode_Float865Output_1113);

ProductNode_Float866: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float866weight,vb3,ProductNode_Float866Output_1114);

ProductNode_Float867: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float867weight,ProductNode_Float7Output_8,ProductNode_Float867Output_1115);

ProductNode_Float868: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float868weight,ProductNode_Float8Output_9,ProductNode_Float868Output_1116);

SumNode_Float248: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float9Output_10,ProductNode_Float6Output_7,SumNode_Float248Output_1117);

ProductNode_Float869: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float1Output_11,ProductNode_Float3Output_4,ProductNode_Float869Output_1118);

ProductNode_Float870: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float870weight,ProductNode_Float10Output_12,ProductNode_Float870Output_1119);

ProductNode_Float871: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float871weight,v8,ProductNode_Float871Output_1120);

ProductNode_Float872: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float872weight,vb8,ProductNode_Float872Output_1121);

SumNode_Float249: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float13Output_15,ProductNode_Float12Output_14,SumNode_Float249Output_1122);

ProductNode_Float873: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb7,SumNode_Float2Output_16,ProductNode_Float873Output_1123);

ProductNode_Float874: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float874weight,v3,ProductNode_Float874Output_1124);

ProductNode_Float875: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float875weight,ProductNode_Float4Output_5,ProductNode_Float875Output_1125);

ProductNode_Float876: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float876weight,ProductNode_Float16Output_19,ProductNode_Float876Output_1126);

ProductNode_Float877: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float877weight,vb3,ProductNode_Float877Output_1127);

ProductNode_Float878: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float878weight,ProductNode_Float7Output_8,ProductNode_Float878Output_1128);

ProductNode_Float879: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float879weight,ProductNode_Float19Output_22,ProductNode_Float879Output_1129);

SumNode_Float250: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float20Output_23,ProductNode_Float17Output_20,SumNode_Float250Output_1130);

ProductNode_Float880: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float3Output_24,ProductNode_Float14Output_17,ProductNode_Float880Output_1131);

ProductNode_Float881: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float881weight,ProductNode_Float21Output_25,ProductNode_Float881Output_1132);

SumNode_Float251: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float595Output_764,ProductNode_Float584Output_751,SumNode_Float251Output_1133);

ProductNode_Float882: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float169Output_765,ProductNode_Float0Output_0,ProductNode_Float882Output_1134);

ProductNode_Float883: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float883weight,ProductNode_Float596Output_766,ProductNode_Float883Output_1135);

ProductNode_Float884: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float884weight,vb4,ProductNode_Float884Output_1136);

ProductNode_Float885: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float885weight,v8,ProductNode_Float885Output_1137);

ProductNode_Float886: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float886weight,vb8,ProductNode_Float886Output_1138);

SumNode_Float252: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float27Output_32,ProductNode_Float26Output_31,SumNode_Float252Output_1139);

ProductNode_Float887: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v7,SumNode_Float5Output_33,ProductNode_Float887Output_1140);

ProductNode_Float888: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float888weight,v3,ProductNode_Float888Output_1141);

ProductNode_Float889: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float889weight,ProductNode_Float29Output_35,ProductNode_Float889Output_1142);

ProductNode_Float890: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float890weight,ProductNode_Float30Output_36,ProductNode_Float890Output_1143);

ProductNode_Float891: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float891weight,vb3,ProductNode_Float891Output_1144);

ProductNode_Float892: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float892weight,ProductNode_Float32Output_38,ProductNode_Float892Output_1145);

ProductNode_Float893: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float893weight,ProductNode_Float33Output_39,ProductNode_Float893Output_1146);

SumNode_Float253: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float34Output_40,ProductNode_Float31Output_37,SumNode_Float253Output_1147);

ProductNode_Float894: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float6Output_41,ProductNode_Float28Output_34,ProductNode_Float894Output_1148);

ProductNode_Float895: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float895weight,ProductNode_Float35Output_42,ProductNode_Float895Output_1149);

ProductNode_Float896: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float896weight,v8,ProductNode_Float896Output_1150);

ProductNode_Float897: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float897weight,vb8,ProductNode_Float897Output_1151);

SumNode_Float254: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float38Output_45,ProductNode_Float37Output_44,SumNode_Float254Output_1152);

ProductNode_Float898: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb7,SumNode_Float7Output_46,ProductNode_Float898Output_1153);

ProductNode_Float899: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float899weight,v3,ProductNode_Float899Output_1154);

ProductNode_Float900: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float900weight,ProductNode_Float29Output_35,ProductNode_Float900Output_1155);

ProductNode_Float901: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float901weight,ProductNode_Float41Output_49,ProductNode_Float901Output_1156);

ProductNode_Float902: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float902weight,vb3,ProductNode_Float902Output_1157);

ProductNode_Float903: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float903weight,ProductNode_Float32Output_38,ProductNode_Float903Output_1158);

ProductNode_Float904: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float904weight,ProductNode_Float44Output_52,ProductNode_Float904Output_1159);

SumNode_Float255: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float45Output_53,ProductNode_Float42Output_50,SumNode_Float255Output_1160);

ProductNode_Float905: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float8Output_54,ProductNode_Float39Output_47,ProductNode_Float905Output_1161);

ProductNode_Float906: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float906weight,ProductNode_Float46Output_55,ProductNode_Float906Output_1162);

SumNode_Float256: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float620Output_794,ProductNode_Float609Output_781,SumNode_Float256Output_1163);

ProductNode_Float907: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float174Output_795,ProductNode_Float25Output_30,ProductNode_Float907Output_1164);

ProductNode_Float908: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float908weight,ProductNode_Float621Output_796,ProductNode_Float908Output_1165);

SumNode_Float257: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float908Output_1165,ProductNode_Float883Output_1135,SumNode_Float257Output_1166);

ProductNode_Float909: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v5,SumNode_Float257Output_1166,ProductNode_Float909Output_1167);

ProductNode_Float910: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float910weight,ProductNode_Float909Output_1167,ProductNode_Float910Output_1168);

ProductNode_Float911: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float911weight,v4,ProductNode_Float911Output_1169);

ProductNode_Float912: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float912weight,v8,ProductNode_Float912Output_1170);

ProductNode_Float913: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float913weight,vb8,ProductNode_Float913Output_1171);

SumNode_Float258: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float54Output_65,ProductNode_Float53Output_64,SumNode_Float258Output_1172);

ProductNode_Float914: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v7,SumNode_Float11Output_66,ProductNode_Float914Output_1173);

ProductNode_Float915: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float915weight,v3,ProductNode_Float915Output_1174);

ProductNode_Float916: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float916weight,ProductNode_Float4Output_5,ProductNode_Float916Output_1175);

ProductNode_Float917: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float917weight,ProductNode_Float5Output_6,ProductNode_Float917Output_1176);

ProductNode_Float918: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float918weight,vb3,ProductNode_Float918Output_1177);

ProductNode_Float919: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float919weight,ProductNode_Float7Output_8,ProductNode_Float919Output_1178);

ProductNode_Float920: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float920weight,ProductNode_Float8Output_9,ProductNode_Float920Output_1179);

SumNode_Float259: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float61Output_73,ProductNode_Float58Output_70,SumNode_Float259Output_1180);

ProductNode_Float921: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float12Output_74,ProductNode_Float55Output_67,ProductNode_Float921Output_1181);

ProductNode_Float922: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float922weight,ProductNode_Float62Output_75,ProductNode_Float922Output_1182);

ProductNode_Float923: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float923weight,v8,ProductNode_Float923Output_1183);

ProductNode_Float924: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float924weight,vb8,ProductNode_Float924Output_1184);

SumNode_Float260: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float65Output_78,ProductNode_Float64Output_77,SumNode_Float260Output_1185);

ProductNode_Float925: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb7,SumNode_Float13Output_79,ProductNode_Float925Output_1186);

ProductNode_Float926: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float926weight,v3,ProductNode_Float926Output_1187);

ProductNode_Float927: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float927weight,ProductNode_Float4Output_5,ProductNode_Float927Output_1188);

ProductNode_Float928: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float928weight,ProductNode_Float16Output_19,ProductNode_Float928Output_1189);

ProductNode_Float929: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float929weight,vb3,ProductNode_Float929Output_1190);

ProductNode_Float930: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float930weight,ProductNode_Float7Output_8,ProductNode_Float930Output_1191);

ProductNode_Float931: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float931weight,ProductNode_Float19Output_22,ProductNode_Float931Output_1192);

SumNode_Float261: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float72Output_86,ProductNode_Float69Output_83,SumNode_Float261Output_1193);

ProductNode_Float932: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float14Output_87,ProductNode_Float66Output_80,ProductNode_Float932Output_1194);

ProductNode_Float933: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float933weight,ProductNode_Float73Output_88,ProductNode_Float933Output_1195);

SumNode_Float262: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float647Output_827,ProductNode_Float636Output_814,SumNode_Float262Output_1196);

ProductNode_Float934: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float180Output_828,ProductNode_Float0Output_0,ProductNode_Float934Output_1197);

ProductNode_Float935: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float935weight,ProductNode_Float648Output_829,ProductNode_Float935Output_1198);

ProductNode_Float936: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float936weight,vb4,ProductNode_Float936Output_1199);

ProductNode_Float937: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float937weight,v8,ProductNode_Float937Output_1200);

ProductNode_Float938: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float938weight,vb8,ProductNode_Float938Output_1201);

SumNode_Float263: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float79Output_95,ProductNode_Float78Output_94,SumNode_Float263Output_1202);

ProductNode_Float939: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v7,SumNode_Float16Output_96,ProductNode_Float939Output_1203);

ProductNode_Float940: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float940weight,v3,ProductNode_Float940Output_1204);

ProductNode_Float941: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float941weight,ProductNode_Float29Output_35,ProductNode_Float941Output_1205);

ProductNode_Float942: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float942weight,ProductNode_Float30Output_36,ProductNode_Float942Output_1206);

ProductNode_Float943: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float943weight,vb3,ProductNode_Float943Output_1207);

ProductNode_Float944: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float944weight,ProductNode_Float32Output_38,ProductNode_Float944Output_1208);

ProductNode_Float945: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float945weight,ProductNode_Float33Output_39,ProductNode_Float945Output_1209);

SumNode_Float264: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float86Output_103,ProductNode_Float83Output_100,SumNode_Float264Output_1210);

ProductNode_Float946: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float17Output_104,ProductNode_Float80Output_97,ProductNode_Float946Output_1211);

ProductNode_Float947: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float947weight,ProductNode_Float87Output_105,ProductNode_Float947Output_1212);

ProductNode_Float948: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float948weight,v8,ProductNode_Float948Output_1213);

ProductNode_Float949: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float949weight,vb8,ProductNode_Float949Output_1214);

SumNode_Float265: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float90Output_108,ProductNode_Float89Output_107,SumNode_Float265Output_1215);

ProductNode_Float950: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb7,SumNode_Float18Output_109,ProductNode_Float950Output_1216);

ProductNode_Float951: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float951weight,v3,ProductNode_Float951Output_1217);

ProductNode_Float952: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float952weight,ProductNode_Float29Output_35,ProductNode_Float952Output_1218);

ProductNode_Float953: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float953weight,ProductNode_Float41Output_49,ProductNode_Float953Output_1219);

ProductNode_Float954: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float954weight,vb3,ProductNode_Float954Output_1220);

ProductNode_Float955: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float955weight,ProductNode_Float32Output_38,ProductNode_Float955Output_1221);

ProductNode_Float956: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float956weight,ProductNode_Float44Output_52,ProductNode_Float956Output_1222);

SumNode_Float266: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float97Output_116,ProductNode_Float94Output_113,SumNode_Float266Output_1223);

ProductNode_Float957: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float19Output_117,ProductNode_Float91Output_110,ProductNode_Float957Output_1224);

ProductNode_Float958: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float958weight,ProductNode_Float98Output_118,ProductNode_Float958Output_1225);

SumNode_Float267: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float672Output_857,ProductNode_Float661Output_844,SumNode_Float267Output_1226);

ProductNode_Float959: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float185Output_858,ProductNode_Float25Output_30,ProductNode_Float959Output_1227);

ProductNode_Float960: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float960weight,ProductNode_Float673Output_859,ProductNode_Float960Output_1228);

SumNode_Float268: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float960Output_1228,ProductNode_Float935Output_1198,SumNode_Float268Output_1229);

ProductNode_Float961: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb5,SumNode_Float268Output_1229,ProductNode_Float961Output_1230);

ProductNode_Float962: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float962weight,ProductNode_Float961Output_1230,ProductNode_Float962Output_1231);

SumNode_Float269: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float962Output_1231,ProductNode_Float910Output_1168,SumNode_Float269Output_1232);

ProductNode_Float963: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb16,SumNode_Float269Output_1232,ProductNode_Float963Output_1233);

ProductNode_Float964: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float964weight,v11,ProductNode_Float964Output_1234);

ProductNode_Float965: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float965weight,vb11,ProductNode_Float965Output_1235);

SumNode_Float270: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float679Output_867,ProductNode_Float678Output_866,SumNode_Float270Output_1236);

ProductNode_Float966: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v12,SumNode_Float188Output_868,ProductNode_Float966Output_1237);

ProductNode_Float967: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float967weight,ProductNode_Float680Output_869,ProductNode_Float967Output_1238);

ProductNode_Float968: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float968weight,v2,ProductNode_Float968Output_1239);

ProductNode_Float969: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float969weight,vb2,ProductNode_Float969Output_1240);

SumNode_Float271: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float110Output_134,ProductNode_Float109Output_133,SumNode_Float271Output_1241);

ProductNode_Float970: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float24Output_135,ProductNode_Float681Output_870,ProductNode_Float970Output_1242);

ProductNode_Float971: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float971weight,v11,ProductNode_Float971Output_1243);

ProductNode_Float972: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float972weight,vb11,ProductNode_Float972Output_1244);

SumNode_Float272: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float686Output_876,ProductNode_Float685Output_875,SumNode_Float272Output_1245);

ProductNode_Float973: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb12,SumNode_Float190Output_877,ProductNode_Float973Output_1246);

ProductNode_Float974: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float974weight,ProductNode_Float687Output_878,ProductNode_Float974Output_1247);

ProductNode_Float975: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float975weight,v2,ProductNode_Float975Output_1248);

ProductNode_Float976: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float976weight,vb2,ProductNode_Float976Output_1249);

SumNode_Float273: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float117Output_143,ProductNode_Float116Output_142,SumNode_Float273Output_1250);

ProductNode_Float977: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float26Output_144,ProductNode_Float688Output_879,ProductNode_Float977Output_1251);

SumNode_Float274: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float691Output_883,ProductNode_Float684Output_874,SumNode_Float274Output_1252);

ProductNode_Float978: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v13,SumNode_Float192Output_884,ProductNode_Float978Output_1253);

ProductNode_Float979: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float979weight,ProductNode_Float692Output_885,ProductNode_Float979Output_1254);

ProductNode_Float980: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float980weight,v11,ProductNode_Float980Output_1255);

ProductNode_Float981: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float981weight,vb11,ProductNode_Float981Output_1256);

SumNode_Float275: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float695Output_888,ProductNode_Float694Output_887,SumNode_Float275Output_1257);

ProductNode_Float982: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v12,SumNode_Float193Output_889,ProductNode_Float982Output_1258);

ProductNode_Float983: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float983weight,ProductNode_Float696Output_890,ProductNode_Float983Output_1259);

ProductNode_Float984: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float984weight,v2,ProductNode_Float984Output_1260);

ProductNode_Float985: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float985weight,vb2,ProductNode_Float985Output_1261);

SumNode_Float276: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float126Output_155,ProductNode_Float125Output_154,SumNode_Float276Output_1262);

ProductNode_Float986: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float29Output_156,ProductNode_Float697Output_891,ProductNode_Float986Output_1263);

ProductNode_Float987: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float987weight,v11,ProductNode_Float987Output_1264);

ProductNode_Float988: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float988weight,vb11,ProductNode_Float988Output_1265);

SumNode_Float277: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float702Output_897,ProductNode_Float701Output_896,SumNode_Float277Output_1266);

ProductNode_Float989: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb12,SumNode_Float195Output_898,ProductNode_Float989Output_1267);

ProductNode_Float990: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float990weight,ProductNode_Float703Output_899,ProductNode_Float990Output_1268);

ProductNode_Float991: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float991weight,v2,ProductNode_Float991Output_1269);

ProductNode_Float992: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float992weight,vb2,ProductNode_Float992Output_1270);

SumNode_Float278: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float133Output_164,ProductNode_Float132Output_163,SumNode_Float278Output_1271);

ProductNode_Float993: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float31Output_165,ProductNode_Float704Output_900,ProductNode_Float993Output_1272);

SumNode_Float279: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float707Output_904,ProductNode_Float700Output_895,SumNode_Float279Output_1273);

ProductNode_Float994: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb13,SumNode_Float197Output_905,ProductNode_Float994Output_1274);

ProductNode_Float995: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float995weight,ProductNode_Float708Output_906,ProductNode_Float995Output_1275);

SumNode_Float280: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float709Output_907,ProductNode_Float693Output_886,SumNode_Float280Output_1276);

ProductNode_Float996: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v10,SumNode_Float198Output_908,ProductNode_Float996Output_1277);

ProductNode_Float997: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float997weight,v1,ProductNode_Float997Output_1278);

ProductNode_Float998: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float998weight,vb1,ProductNode_Float998Output_1279);

SumNode_Float281: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float139Output_173,ProductNode_Float138Output_172,SumNode_Float281Output_1280);

ProductNode_Float999: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v9,SumNode_Float34Output_174,ProductNode_Float999Output_1281);

ProductNode_Float1000: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1000weight,ProductNode_Float140Output_175,ProductNode_Float1000Output_1282);

ProductNode_Float1001: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1001weight,ProductNode_Float141Output_176,ProductNode_Float1001Output_1283);

ProductNode_Float1002: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1002weight,v1,ProductNode_Float1002Output_1284);

ProductNode_Float1003: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1003weight,vb1,ProductNode_Float1003Output_1285);

SumNode_Float282: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float144Output_179,ProductNode_Float143Output_178,SumNode_Float282Output_1286);

ProductNode_Float1004: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb9,SumNode_Float35Output_180,ProductNode_Float1004Output_1287);

ProductNode_Float1005: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1005weight,ProductNode_Float145Output_181,ProductNode_Float1005Output_1288);

ProductNode_Float1006: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1006weight,ProductNode_Float146Output_182,ProductNode_Float1006Output_1289);

SumNode_Float283: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float147Output_183,ProductNode_Float142Output_177,SumNode_Float283Output_1290);

ProductNode_Float1007: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float36Output_184,ProductNode_Float710Output_909,ProductNode_Float1007Output_1291);

ProductNode_Float1008: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1008weight,v11,ProductNode_Float1008Output_1292);

ProductNode_Float1009: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1009weight,vb11,ProductNode_Float1009Output_1293);

SumNode_Float284: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float679Output_867,ProductNode_Float678Output_866,SumNode_Float284Output_1294);

ProductNode_Float1010: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v12,SumNode_Float188Output_868,ProductNode_Float1010Output_1295);

ProductNode_Float1011: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1011weight,ProductNode_Float680Output_869,ProductNode_Float1011Output_1296);

ProductNode_Float1012: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1012weight,v2,ProductNode_Float1012Output_1297);

ProductNode_Float1013: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1013weight,vb2,ProductNode_Float1013Output_1298);

SumNode_Float285: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float110Output_134,ProductNode_Float109Output_133,SumNode_Float285Output_1299);

ProductNode_Float1014: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float24Output_135,ProductNode_Float681Output_870,ProductNode_Float1014Output_1300);

ProductNode_Float1015: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1015weight,v11,ProductNode_Float1015Output_1301);

ProductNode_Float1016: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1016weight,vb11,ProductNode_Float1016Output_1302);

SumNode_Float286: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float686Output_876,ProductNode_Float685Output_875,SumNode_Float286Output_1303);

ProductNode_Float1017: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb12,SumNode_Float190Output_877,ProductNode_Float1017Output_1304);

ProductNode_Float1018: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1018weight,ProductNode_Float687Output_878,ProductNode_Float1018Output_1305);

ProductNode_Float1019: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1019weight,v2,ProductNode_Float1019Output_1306);

ProductNode_Float1020: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1020weight,vb2,ProductNode_Float1020Output_1307);

SumNode_Float287: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float117Output_143,ProductNode_Float116Output_142,SumNode_Float287Output_1308);

ProductNode_Float1021: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float26Output_144,ProductNode_Float688Output_879,ProductNode_Float1021Output_1309);

SumNode_Float288: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float691Output_883,ProductNode_Float684Output_874,SumNode_Float288Output_1310);

ProductNode_Float1022: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v13,SumNode_Float192Output_884,ProductNode_Float1022Output_1311);

ProductNode_Float1023: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1023weight,ProductNode_Float692Output_885,ProductNode_Float1023Output_1312);

ProductNode_Float1024: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1024weight,v11,ProductNode_Float1024Output_1313);

ProductNode_Float1025: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1025weight,vb11,ProductNode_Float1025Output_1314);

SumNode_Float289: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float695Output_888,ProductNode_Float694Output_887,SumNode_Float289Output_1315);

ProductNode_Float1026: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v12,SumNode_Float193Output_889,ProductNode_Float1026Output_1316);

ProductNode_Float1027: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1027weight,ProductNode_Float696Output_890,ProductNode_Float1027Output_1317);

ProductNode_Float1028: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1028weight,v2,ProductNode_Float1028Output_1318);

ProductNode_Float1029: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1029weight,vb2,ProductNode_Float1029Output_1319);

SumNode_Float290: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float126Output_155,ProductNode_Float125Output_154,SumNode_Float290Output_1320);

ProductNode_Float1030: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float29Output_156,ProductNode_Float697Output_891,ProductNode_Float1030Output_1321);

ProductNode_Float1031: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1031weight,v11,ProductNode_Float1031Output_1322);

ProductNode_Float1032: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1032weight,vb11,ProductNode_Float1032Output_1323);

SumNode_Float291: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float702Output_897,ProductNode_Float701Output_896,SumNode_Float291Output_1324);

ProductNode_Float1033: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb12,SumNode_Float195Output_898,ProductNode_Float1033Output_1325);

ProductNode_Float1034: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1034weight,ProductNode_Float703Output_899,ProductNode_Float1034Output_1326);

ProductNode_Float1035: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1035weight,v2,ProductNode_Float1035Output_1327);

ProductNode_Float1036: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1036weight,vb2,ProductNode_Float1036Output_1328);

SumNode_Float292: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float133Output_164,ProductNode_Float132Output_163,SumNode_Float292Output_1329);

ProductNode_Float1037: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float31Output_165,ProductNode_Float704Output_900,ProductNode_Float1037Output_1330);

SumNode_Float293: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float707Output_904,ProductNode_Float700Output_895,SumNode_Float293Output_1331);

ProductNode_Float1038: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb13,SumNode_Float197Output_905,ProductNode_Float1038Output_1332);

ProductNode_Float1039: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1039weight,ProductNode_Float708Output_906,ProductNode_Float1039Output_1333);

SumNode_Float294: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float753Output_965,ProductNode_Float737Output_944,SumNode_Float294Output_1334);

ProductNode_Float1040: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb10,SumNode_Float212Output_966,ProductNode_Float1040Output_1335);

ProductNode_Float1041: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1041weight,v1,ProductNode_Float1041Output_1336);

ProductNode_Float1042: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1042weight,vb1,ProductNode_Float1042Output_1337);

SumNode_Float295: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float183Output_231,ProductNode_Float182Output_230,SumNode_Float295Output_1338);

ProductNode_Float1043: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v9,SumNode_Float48Output_232,ProductNode_Float1043Output_1339);

ProductNode_Float1044: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1044weight,ProductNode_Float184Output_233,ProductNode_Float1044Output_1340);

ProductNode_Float1045: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1045weight,ProductNode_Float185Output_234,ProductNode_Float1045Output_1341);

ProductNode_Float1046: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1046weight,v1,ProductNode_Float1046Output_1342);

ProductNode_Float1047: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1047weight,vb1,ProductNode_Float1047Output_1343);

SumNode_Float296: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float188Output_237,ProductNode_Float187Output_236,SumNode_Float296Output_1344);

ProductNode_Float1048: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb9,SumNode_Float49Output_238,ProductNode_Float1048Output_1345);

ProductNode_Float1049: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1049weight,ProductNode_Float189Output_239,ProductNode_Float1049Output_1346);

ProductNode_Float1050: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1050weight,ProductNode_Float190Output_240,ProductNode_Float1050Output_1347);

SumNode_Float297: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float191Output_241,ProductNode_Float186Output_235,SumNode_Float297Output_1348);

ProductNode_Float1051: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float50Output_242,ProductNode_Float754Output_967,ProductNode_Float1051Output_1349);

SumNode_Float298: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float765Output_981,ProductNode_Float721Output_923,SumNode_Float298Output_1350);

ProductNode_Float1052: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v15,SumNode_Float216Output_982,ProductNode_Float1052Output_1351);

ProductNode_Float1053: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1053weight,ProductNode_Float766Output_983,ProductNode_Float1053Output_1352);

ProductNode_Float1054: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1054weight,v11,ProductNode_Float1054Output_1353);

ProductNode_Float1055: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1055weight,vb11,ProductNode_Float1055Output_1354);

SumNode_Float299: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float679Output_867,ProductNode_Float678Output_866,SumNode_Float299Output_1355);

ProductNode_Float1056: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v12,SumNode_Float188Output_868,ProductNode_Float1056Output_1356);

ProductNode_Float1057: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1057weight,ProductNode_Float680Output_869,ProductNode_Float1057Output_1357);

ProductNode_Float1058: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1058weight,v2,ProductNode_Float1058Output_1358);

ProductNode_Float1059: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1059weight,vb2,ProductNode_Float1059Output_1359);

SumNode_Float300: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float200Output_253,ProductNode_Float199Output_252,SumNode_Float300Output_1360);

ProductNode_Float1060: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float53Output_254,ProductNode_Float681Output_870,ProductNode_Float1060Output_1361);

ProductNode_Float1061: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1061weight,v11,ProductNode_Float1061Output_1362);

ProductNode_Float1062: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1062weight,vb11,ProductNode_Float1062Output_1363);

SumNode_Float301: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float686Output_876,ProductNode_Float685Output_875,SumNode_Float301Output_1364);

ProductNode_Float1063: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb12,SumNode_Float190Output_877,ProductNode_Float1063Output_1365);

ProductNode_Float1064: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1064weight,ProductNode_Float687Output_878,ProductNode_Float1064Output_1366);

ProductNode_Float1065: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1065weight,v2,ProductNode_Float1065Output_1367);

ProductNode_Float1066: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1066weight,vb2,ProductNode_Float1066Output_1368);

SumNode_Float302: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float207Output_262,ProductNode_Float206Output_261,SumNode_Float302Output_1369);

ProductNode_Float1067: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float55Output_263,ProductNode_Float688Output_879,ProductNode_Float1067Output_1370);

SumNode_Float303: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float781Output_1002,ProductNode_Float774Output_993,SumNode_Float303Output_1371);

ProductNode_Float1068: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v13,SumNode_Float221Output_1003,ProductNode_Float1068Output_1372);

ProductNode_Float1069: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1069weight,ProductNode_Float782Output_1004,ProductNode_Float1069Output_1373);

ProductNode_Float1070: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1070weight,v11,ProductNode_Float1070Output_1374);

ProductNode_Float1071: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1071weight,vb11,ProductNode_Float1071Output_1375);

SumNode_Float304: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float695Output_888,ProductNode_Float694Output_887,SumNode_Float304Output_1376);

ProductNode_Float1072: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v12,SumNode_Float193Output_889,ProductNode_Float1072Output_1377);

ProductNode_Float1073: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1073weight,ProductNode_Float696Output_890,ProductNode_Float1073Output_1378);

ProductNode_Float1074: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1074weight,v2,ProductNode_Float1074Output_1379);

ProductNode_Float1075: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1075weight,vb2,ProductNode_Float1075Output_1380);

SumNode_Float305: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float216Output_274,ProductNode_Float215Output_273,SumNode_Float305Output_1381);

ProductNode_Float1076: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float58Output_275,ProductNode_Float697Output_891,ProductNode_Float1076Output_1382);

ProductNode_Float1077: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1077weight,v11,ProductNode_Float1077Output_1383);

ProductNode_Float1078: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1078weight,vb11,ProductNode_Float1078Output_1384);

SumNode_Float306: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float702Output_897,ProductNode_Float701Output_896,SumNode_Float306Output_1385);

ProductNode_Float1079: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb12,SumNode_Float195Output_898,ProductNode_Float1079Output_1386);

ProductNode_Float1080: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1080weight,ProductNode_Float703Output_899,ProductNode_Float1080Output_1387);

ProductNode_Float1081: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1081weight,v2,ProductNode_Float1081Output_1388);

ProductNode_Float1082: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1082weight,vb2,ProductNode_Float1082Output_1389);

SumNode_Float307: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float223Output_283,ProductNode_Float222Output_282,SumNode_Float307Output_1390);

ProductNode_Float1083: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float60Output_284,ProductNode_Float704Output_900,ProductNode_Float1083Output_1391);

SumNode_Float308: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float797Output_1023,ProductNode_Float790Output_1014,SumNode_Float308Output_1392);

ProductNode_Float1084: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb13,SumNode_Float226Output_1024,ProductNode_Float1084Output_1393);

ProductNode_Float1085: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1085weight,ProductNode_Float798Output_1025,ProductNode_Float1085Output_1394);

SumNode_Float309: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float799Output_1026,ProductNode_Float783Output_1005,SumNode_Float309Output_1395);

ProductNode_Float1086: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v10,SumNode_Float227Output_1027,ProductNode_Float1086Output_1396);

ProductNode_Float1087: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1087weight,v1,ProductNode_Float1087Output_1397);

ProductNode_Float1088: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1088weight,vb1,ProductNode_Float1088Output_1398);

SumNode_Float310: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float139Output_173,ProductNode_Float138Output_172,SumNode_Float310Output_1399);

ProductNode_Float1089: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v9,SumNode_Float34Output_174,ProductNode_Float1089Output_1400);

ProductNode_Float1090: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1090weight,ProductNode_Float140Output_175,ProductNode_Float1090Output_1401);

ProductNode_Float1091: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1091weight,ProductNode_Float231Output_295,ProductNode_Float1091Output_1402);

ProductNode_Float1092: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1092weight,v1,ProductNode_Float1092Output_1403);

ProductNode_Float1093: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1093weight,vb1,ProductNode_Float1093Output_1404);

SumNode_Float311: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float144Output_179,ProductNode_Float143Output_178,SumNode_Float311Output_1405);

ProductNode_Float1094: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb9,SumNode_Float35Output_180,ProductNode_Float1094Output_1406);

ProductNode_Float1095: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1095weight,ProductNode_Float145Output_181,ProductNode_Float1095Output_1407);

ProductNode_Float1096: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1096weight,ProductNode_Float236Output_301,ProductNode_Float1096Output_1408);

SumNode_Float312: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float237Output_302,ProductNode_Float232Output_296,SumNode_Float312Output_1409);

ProductNode_Float1097: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float65Output_303,ProductNode_Float800Output_1028,ProductNode_Float1097Output_1410);

ProductNode_Float1098: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1098weight,v11,ProductNode_Float1098Output_1411);

ProductNode_Float1099: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1099weight,vb11,ProductNode_Float1099Output_1412);

SumNode_Float313: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float679Output_867,ProductNode_Float678Output_866,SumNode_Float313Output_1413);

ProductNode_Float1100: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v12,SumNode_Float188Output_868,ProductNode_Float1100Output_1414);

ProductNode_Float1101: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1101weight,ProductNode_Float680Output_869,ProductNode_Float1101Output_1415);

ProductNode_Float1102: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1102weight,v2,ProductNode_Float1102Output_1416);

ProductNode_Float1103: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1103weight,vb2,ProductNode_Float1103Output_1417);

SumNode_Float314: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float200Output_253,ProductNode_Float199Output_252,SumNode_Float314Output_1418);

ProductNode_Float1104: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float53Output_254,ProductNode_Float681Output_870,ProductNode_Float1104Output_1419);

ProductNode_Float1105: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1105weight,v11,ProductNode_Float1105Output_1420);

ProductNode_Float1106: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1106weight,vb11,ProductNode_Float1106Output_1421);

SumNode_Float315: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float686Output_876,ProductNode_Float685Output_875,SumNode_Float315Output_1422);

ProductNode_Float1107: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb12,SumNode_Float190Output_877,ProductNode_Float1107Output_1423);

ProductNode_Float1108: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1108weight,ProductNode_Float687Output_878,ProductNode_Float1108Output_1424);

ProductNode_Float1109: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1109weight,v2,ProductNode_Float1109Output_1425);

ProductNode_Float1110: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1110weight,vb2,ProductNode_Float1110Output_1426);

SumNode_Float316: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float207Output_262,ProductNode_Float206Output_261,SumNode_Float316Output_1427);

ProductNode_Float1111: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float55Output_263,ProductNode_Float688Output_879,ProductNode_Float1111Output_1428);

SumNode_Float317: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float781Output_1002,ProductNode_Float774Output_993,SumNode_Float317Output_1429);

ProductNode_Float1112: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v13,SumNode_Float221Output_1003,ProductNode_Float1112Output_1430);

ProductNode_Float1113: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1113weight,ProductNode_Float782Output_1004,ProductNode_Float1113Output_1431);

ProductNode_Float1114: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1114weight,v11,ProductNode_Float1114Output_1432);

ProductNode_Float1115: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1115weight,vb11,ProductNode_Float1115Output_1433);

SumNode_Float318: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float695Output_888,ProductNode_Float694Output_887,SumNode_Float318Output_1434);

ProductNode_Float1116: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v12,SumNode_Float193Output_889,ProductNode_Float1116Output_1435);

ProductNode_Float1117: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1117weight,ProductNode_Float696Output_890,ProductNode_Float1117Output_1436);

ProductNode_Float1118: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1118weight,v2,ProductNode_Float1118Output_1437);

ProductNode_Float1119: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1119weight,vb2,ProductNode_Float1119Output_1438);

SumNode_Float319: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float216Output_274,ProductNode_Float215Output_273,SumNode_Float319Output_1439);

ProductNode_Float1120: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float58Output_275,ProductNode_Float697Output_891,ProductNode_Float1120Output_1440);

ProductNode_Float1121: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1121weight,v11,ProductNode_Float1121Output_1441);

ProductNode_Float1122: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1122weight,vb11,ProductNode_Float1122Output_1442);

SumNode_Float320: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float702Output_897,ProductNode_Float701Output_896,SumNode_Float320Output_1443);

ProductNode_Float1123: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb12,SumNode_Float195Output_898,ProductNode_Float1123Output_1444);

ProductNode_Float1124: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1124weight,ProductNode_Float703Output_899,ProductNode_Float1124Output_1445);

ProductNode_Float1125: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1125weight,v2,ProductNode_Float1125Output_1446);

ProductNode_Float1126: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1126weight,vb2,ProductNode_Float1126Output_1447);

SumNode_Float321: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float223Output_283,ProductNode_Float222Output_282,SumNode_Float321Output_1448);

ProductNode_Float1127: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float60Output_284,ProductNode_Float704Output_900,ProductNode_Float1127Output_1449);

SumNode_Float322: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float797Output_1023,ProductNode_Float790Output_1014,SumNode_Float322Output_1450);

ProductNode_Float1128: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb13,SumNode_Float226Output_1024,ProductNode_Float1128Output_1451);

ProductNode_Float1129: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1129weight,ProductNode_Float798Output_1025,ProductNode_Float1129Output_1452);

SumNode_Float323: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float843Output_1084,ProductNode_Float827Output_1063,SumNode_Float323Output_1453);

ProductNode_Float1130: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb10,SumNode_Float241Output_1085,ProductNode_Float1130Output_1454);

ProductNode_Float1131: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1131weight,v1,ProductNode_Float1131Output_1455);

ProductNode_Float1132: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1132weight,vb1,ProductNode_Float1132Output_1456);

SumNode_Float324: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float183Output_231,ProductNode_Float182Output_230,SumNode_Float324Output_1457);

ProductNode_Float1133: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v9,SumNode_Float48Output_232,ProductNode_Float1133Output_1458);

ProductNode_Float1134: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1134weight,ProductNode_Float184Output_233,ProductNode_Float1134Output_1459);

ProductNode_Float1135: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1135weight,ProductNode_Float275Output_353,ProductNode_Float1135Output_1460);

ProductNode_Float1136: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1136weight,v1,ProductNode_Float1136Output_1461);

ProductNode_Float1137: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1137weight,vb1,ProductNode_Float1137Output_1462);

SumNode_Float325: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float188Output_237,ProductNode_Float187Output_236,SumNode_Float325Output_1463);

ProductNode_Float1138: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb9,SumNode_Float49Output_238,ProductNode_Float1138Output_1464);

ProductNode_Float1139: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1139weight,ProductNode_Float189Output_239,ProductNode_Float1139Output_1465);

ProductNode_Float1140: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1140weight,ProductNode_Float280Output_359,ProductNode_Float1140Output_1466);

SumNode_Float326: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float281Output_360,ProductNode_Float276Output_354,SumNode_Float326Output_1467);

ProductNode_Float1141: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float79Output_361,ProductNode_Float844Output_1086,ProductNode_Float1141Output_1468);

SumNode_Float327: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float855Output_1100,ProductNode_Float811Output_1042,SumNode_Float327Output_1469);

ProductNode_Float1142: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb15,SumNode_Float245Output_1101,ProductNode_Float1142Output_1470);

ProductNode_Float1143: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1143weight,ProductNode_Float856Output_1102,ProductNode_Float1143Output_1471);

SumNode_Float328: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1143Output_1471,ProductNode_Float1053Output_1352,SumNode_Float328Output_1472);

ProductNode_Float1144: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float328Output_1472,ProductNode_Float963Output_1233,ProductNode_Float1144Output_1473);

SumNode_Float329: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1144Output_1473,ProductNode_Float858Output_1105,SumNode_Float329Output_1474);

ProductNode_Float1145: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb6,SumNode_Float329Output_1474,ProductNode_Float1145Output_1475);

SumNode_Float330: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1145Output_1475,ProductNode_Float572Output_737,SumNode_Float330Output_1476);

ProductNode_Float1146: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v14,SumNode_Float330Output_1476,ProductNode_Float1146Output_1477);

ProductNode_Float1147: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1147weight,v4,ProductNode_Float1147Output_1478);

ProductNode_Float1148: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1148weight,v8,ProductNode_Float1148Output_1479);

ProductNode_Float1149: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1149weight,vb8,ProductNode_Float1149Output_1480);

SumNode_Float331: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2Output_2,ProductNode_Float1Output_1,SumNode_Float331Output_1481);

ProductNode_Float1150: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v7,SumNode_Float0Output_3,ProductNode_Float1150Output_1482);

ProductNode_Float1151: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1151weight,v3,ProductNode_Float1151Output_1483);

ProductNode_Float1152: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1152weight,ProductNode_Float4Output_5,ProductNode_Float1152Output_1484);

ProductNode_Float1153: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1153weight,ProductNode_Float5Output_6,ProductNode_Float1153Output_1485);

ProductNode_Float1154: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1154weight,vb3,ProductNode_Float1154Output_1486);

ProductNode_Float1155: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1155weight,ProductNode_Float7Output_8,ProductNode_Float1155Output_1487);

ProductNode_Float1156: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1156weight,ProductNode_Float8Output_9,ProductNode_Float1156Output_1488);

SumNode_Float332: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float9Output_10,ProductNode_Float6Output_7,SumNode_Float332Output_1489);

ProductNode_Float1157: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float1Output_11,ProductNode_Float3Output_4,ProductNode_Float1157Output_1490);

ProductNode_Float1158: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1158weight,ProductNode_Float10Output_12,ProductNode_Float1158Output_1491);

ProductNode_Float1159: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1159weight,v8,ProductNode_Float1159Output_1492);

ProductNode_Float1160: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1160weight,vb8,ProductNode_Float1160Output_1493);

SumNode_Float333: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float13Output_15,ProductNode_Float12Output_14,SumNode_Float333Output_1494);

ProductNode_Float1161: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb7,SumNode_Float2Output_16,ProductNode_Float1161Output_1495);

ProductNode_Float1162: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1162weight,v3,ProductNode_Float1162Output_1496);

ProductNode_Float1163: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1163weight,ProductNode_Float4Output_5,ProductNode_Float1163Output_1497);

ProductNode_Float1164: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1164weight,ProductNode_Float16Output_19,ProductNode_Float1164Output_1498);

ProductNode_Float1165: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1165weight,vb3,ProductNode_Float1165Output_1499);

ProductNode_Float1166: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1166weight,ProductNode_Float7Output_8,ProductNode_Float1166Output_1500);

ProductNode_Float1167: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1167weight,ProductNode_Float19Output_22,ProductNode_Float1167Output_1501);

SumNode_Float334: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float20Output_23,ProductNode_Float17Output_20,SumNode_Float334Output_1502);

ProductNode_Float1168: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float3Output_24,ProductNode_Float14Output_17,ProductNode_Float1168Output_1503);

ProductNode_Float1169: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1169weight,ProductNode_Float21Output_25,ProductNode_Float1169Output_1504);

SumNode_Float335: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float22Output_26,ProductNode_Float11Output_13,SumNode_Float335Output_1505);

ProductNode_Float1170: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float4Output_27,ProductNode_Float0Output_0,ProductNode_Float1170Output_1506);

ProductNode_Float1171: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1171weight,ProductNode_Float23Output_28,ProductNode_Float1171Output_1507);

ProductNode_Float1172: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1172weight,vb4,ProductNode_Float1172Output_1508);

ProductNode_Float1173: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1173weight,v8,ProductNode_Float1173Output_1509);

ProductNode_Float1174: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1174weight,vb8,ProductNode_Float1174Output_1510);

SumNode_Float336: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float27Output_32,ProductNode_Float26Output_31,SumNode_Float336Output_1511);

ProductNode_Float1175: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v7,SumNode_Float5Output_33,ProductNode_Float1175Output_1512);

ProductNode_Float1176: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1176weight,v3,ProductNode_Float1176Output_1513);

ProductNode_Float1177: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1177weight,ProductNode_Float29Output_35,ProductNode_Float1177Output_1514);

ProductNode_Float1178: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1178weight,ProductNode_Float30Output_36,ProductNode_Float1178Output_1515);

ProductNode_Float1179: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1179weight,vb3,ProductNode_Float1179Output_1516);

ProductNode_Float1180: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1180weight,ProductNode_Float32Output_38,ProductNode_Float1180Output_1517);

ProductNode_Float1181: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1181weight,ProductNode_Float33Output_39,ProductNode_Float1181Output_1518);

SumNode_Float337: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float34Output_40,ProductNode_Float31Output_37,SumNode_Float337Output_1519);

ProductNode_Float1182: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float6Output_41,ProductNode_Float28Output_34,ProductNode_Float1182Output_1520);

ProductNode_Float1183: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1183weight,ProductNode_Float35Output_42,ProductNode_Float1183Output_1521);

ProductNode_Float1184: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1184weight,v8,ProductNode_Float1184Output_1522);

ProductNode_Float1185: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1185weight,vb8,ProductNode_Float1185Output_1523);

SumNode_Float338: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float38Output_45,ProductNode_Float37Output_44,SumNode_Float338Output_1524);

ProductNode_Float1186: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb7,SumNode_Float7Output_46,ProductNode_Float1186Output_1525);

ProductNode_Float1187: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1187weight,v3,ProductNode_Float1187Output_1526);

ProductNode_Float1188: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1188weight,ProductNode_Float29Output_35,ProductNode_Float1188Output_1527);

ProductNode_Float1189: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1189weight,ProductNode_Float41Output_49,ProductNode_Float1189Output_1528);

ProductNode_Float1190: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1190weight,vb3,ProductNode_Float1190Output_1529);

ProductNode_Float1191: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1191weight,ProductNode_Float32Output_38,ProductNode_Float1191Output_1530);

ProductNode_Float1192: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1192weight,ProductNode_Float44Output_52,ProductNode_Float1192Output_1531);

SumNode_Float339: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float45Output_53,ProductNode_Float42Output_50,SumNode_Float339Output_1532);

ProductNode_Float1193: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float8Output_54,ProductNode_Float39Output_47,ProductNode_Float1193Output_1533);

ProductNode_Float1194: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1194weight,ProductNode_Float46Output_55,ProductNode_Float1194Output_1534);

SumNode_Float340: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float47Output_56,ProductNode_Float36Output_43,SumNode_Float340Output_1535);

ProductNode_Float1195: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float9Output_57,ProductNode_Float25Output_30,ProductNode_Float1195Output_1536);

ProductNode_Float1196: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1196weight,ProductNode_Float48Output_58,ProductNode_Float1196Output_1537);

SumNode_Float341: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float49Output_59,ProductNode_Float24Output_29,SumNode_Float341Output_1538);

ProductNode_Float1197: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v5,SumNode_Float10Output_60,ProductNode_Float1197Output_1539);

ProductNode_Float1198: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1198weight,ProductNode_Float50Output_61,ProductNode_Float1198Output_1540);

ProductNode_Float1199: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1199weight,v4,ProductNode_Float1199Output_1541);

ProductNode_Float1200: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1200weight,v8,ProductNode_Float1200Output_1542);

ProductNode_Float1201: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1201weight,vb8,ProductNode_Float1201Output_1543);

SumNode_Float342: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float54Output_65,ProductNode_Float53Output_64,SumNode_Float342Output_1544);

ProductNode_Float1202: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v7,SumNode_Float11Output_66,ProductNode_Float1202Output_1545);

ProductNode_Float1203: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1203weight,v3,ProductNode_Float1203Output_1546);

ProductNode_Float1204: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1204weight,ProductNode_Float4Output_5,ProductNode_Float1204Output_1547);

ProductNode_Float1205: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1205weight,ProductNode_Float5Output_6,ProductNode_Float1205Output_1548);

ProductNode_Float1206: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1206weight,vb3,ProductNode_Float1206Output_1549);

ProductNode_Float1207: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1207weight,ProductNode_Float7Output_8,ProductNode_Float1207Output_1550);

ProductNode_Float1208: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1208weight,ProductNode_Float8Output_9,ProductNode_Float1208Output_1551);

SumNode_Float343: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float61Output_73,ProductNode_Float58Output_70,SumNode_Float343Output_1552);

ProductNode_Float1209: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float12Output_74,ProductNode_Float55Output_67,ProductNode_Float1209Output_1553);

ProductNode_Float1210: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1210weight,ProductNode_Float62Output_75,ProductNode_Float1210Output_1554);

ProductNode_Float1211: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1211weight,v8,ProductNode_Float1211Output_1555);

ProductNode_Float1212: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1212weight,vb8,ProductNode_Float1212Output_1556);

SumNode_Float344: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float65Output_78,ProductNode_Float64Output_77,SumNode_Float344Output_1557);

ProductNode_Float1213: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb7,SumNode_Float13Output_79,ProductNode_Float1213Output_1558);

ProductNode_Float1214: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1214weight,v3,ProductNode_Float1214Output_1559);

ProductNode_Float1215: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1215weight,ProductNode_Float4Output_5,ProductNode_Float1215Output_1560);

ProductNode_Float1216: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1216weight,ProductNode_Float16Output_19,ProductNode_Float1216Output_1561);

ProductNode_Float1217: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1217weight,vb3,ProductNode_Float1217Output_1562);

ProductNode_Float1218: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1218weight,ProductNode_Float7Output_8,ProductNode_Float1218Output_1563);

ProductNode_Float1219: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1219weight,ProductNode_Float19Output_22,ProductNode_Float1219Output_1564);

SumNode_Float345: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float72Output_86,ProductNode_Float69Output_83,SumNode_Float345Output_1565);

ProductNode_Float1220: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float14Output_87,ProductNode_Float66Output_80,ProductNode_Float1220Output_1566);

ProductNode_Float1221: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1221weight,ProductNode_Float73Output_88,ProductNode_Float1221Output_1567);

SumNode_Float346: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float74Output_89,ProductNode_Float63Output_76,SumNode_Float346Output_1568);

ProductNode_Float1222: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float15Output_90,ProductNode_Float0Output_0,ProductNode_Float1222Output_1569);

ProductNode_Float1223: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1223weight,ProductNode_Float75Output_91,ProductNode_Float1223Output_1570);

ProductNode_Float1224: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1224weight,vb4,ProductNode_Float1224Output_1571);

ProductNode_Float1225: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1225weight,v8,ProductNode_Float1225Output_1572);

ProductNode_Float1226: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1226weight,vb8,ProductNode_Float1226Output_1573);

SumNode_Float347: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float79Output_95,ProductNode_Float78Output_94,SumNode_Float347Output_1574);

ProductNode_Float1227: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v7,SumNode_Float16Output_96,ProductNode_Float1227Output_1575);

ProductNode_Float1228: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1228weight,v3,ProductNode_Float1228Output_1576);

ProductNode_Float1229: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1229weight,ProductNode_Float29Output_35,ProductNode_Float1229Output_1577);

ProductNode_Float1230: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1230weight,ProductNode_Float30Output_36,ProductNode_Float1230Output_1578);

ProductNode_Float1231: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1231weight,vb3,ProductNode_Float1231Output_1579);

ProductNode_Float1232: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1232weight,ProductNode_Float32Output_38,ProductNode_Float1232Output_1580);

ProductNode_Float1233: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1233weight,ProductNode_Float33Output_39,ProductNode_Float1233Output_1581);

SumNode_Float348: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float86Output_103,ProductNode_Float83Output_100,SumNode_Float348Output_1582);

ProductNode_Float1234: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float17Output_104,ProductNode_Float80Output_97,ProductNode_Float1234Output_1583);

ProductNode_Float1235: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1235weight,ProductNode_Float87Output_105,ProductNode_Float1235Output_1584);

ProductNode_Float1236: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1236weight,v8,ProductNode_Float1236Output_1585);

ProductNode_Float1237: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1237weight,vb8,ProductNode_Float1237Output_1586);

SumNode_Float349: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float90Output_108,ProductNode_Float89Output_107,SumNode_Float349Output_1587);

ProductNode_Float1238: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb7,SumNode_Float18Output_109,ProductNode_Float1238Output_1588);

ProductNode_Float1239: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1239weight,v3,ProductNode_Float1239Output_1589);

ProductNode_Float1240: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1240weight,ProductNode_Float29Output_35,ProductNode_Float1240Output_1590);

ProductNode_Float1241: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1241weight,ProductNode_Float41Output_49,ProductNode_Float1241Output_1591);

ProductNode_Float1242: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1242weight,vb3,ProductNode_Float1242Output_1592);

ProductNode_Float1243: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1243weight,ProductNode_Float32Output_38,ProductNode_Float1243Output_1593);

ProductNode_Float1244: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1244weight,ProductNode_Float44Output_52,ProductNode_Float1244Output_1594);

SumNode_Float350: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float97Output_116,ProductNode_Float94Output_113,SumNode_Float350Output_1595);

ProductNode_Float1245: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float19Output_117,ProductNode_Float91Output_110,ProductNode_Float1245Output_1596);

ProductNode_Float1246: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1246weight,ProductNode_Float98Output_118,ProductNode_Float1246Output_1597);

SumNode_Float351: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float99Output_119,ProductNode_Float88Output_106,SumNode_Float351Output_1598);

ProductNode_Float1247: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float20Output_120,ProductNode_Float25Output_30,ProductNode_Float1247Output_1599);

ProductNode_Float1248: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1248weight,ProductNode_Float100Output_121,ProductNode_Float1248Output_1600);

SumNode_Float352: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float101Output_122,ProductNode_Float76Output_92,SumNode_Float352Output_1601);

ProductNode_Float1249: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb5,SumNode_Float21Output_123,ProductNode_Float1249Output_1602);

ProductNode_Float1250: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1250weight,ProductNode_Float102Output_124,ProductNode_Float1250Output_1603);

SumNode_Float353: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1250Output_1603,ProductNode_Float1198Output_1540,SumNode_Float353Output_1604);

ProductNode_Float1251: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v16,SumNode_Float353Output_1604,ProductNode_Float1251Output_1605);

ProductNode_Float1252: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1252weight,v11,ProductNode_Float1252Output_1606);

ProductNode_Float1253: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1253weight,vb11,ProductNode_Float1253Output_1607);

SumNode_Float354: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float106Output_129,ProductNode_Float105Output_128,SumNode_Float354Output_1608);

ProductNode_Float1254: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v12,SumNode_Float23Output_130,ProductNode_Float1254Output_1609);

ProductNode_Float1255: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1255weight,ProductNode_Float107Output_131,ProductNode_Float1255Output_1610);

ProductNode_Float1256: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1256weight,v2,ProductNode_Float1256Output_1611);

ProductNode_Float1257: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1257weight,vb2,ProductNode_Float1257Output_1612);

SumNode_Float355: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float110Output_134,ProductNode_Float109Output_133,SumNode_Float355Output_1613);

ProductNode_Float1258: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float24Output_135,ProductNode_Float108Output_132,ProductNode_Float1258Output_1614);

ProductNode_Float1259: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1259weight,v11,ProductNode_Float1259Output_1615);

ProductNode_Float1260: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1260weight,vb11,ProductNode_Float1260Output_1616);

SumNode_Float356: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float113Output_138,ProductNode_Float112Output_137,SumNode_Float356Output_1617);

ProductNode_Float1261: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb12,SumNode_Float25Output_139,ProductNode_Float1261Output_1618);

ProductNode_Float1262: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1262weight,ProductNode_Float114Output_140,ProductNode_Float1262Output_1619);

ProductNode_Float1263: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1263weight,v2,ProductNode_Float1263Output_1620);

ProductNode_Float1264: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1264weight,vb2,ProductNode_Float1264Output_1621);

SumNode_Float357: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float117Output_143,ProductNode_Float116Output_142,SumNode_Float357Output_1622);

ProductNode_Float1265: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float26Output_144,ProductNode_Float115Output_141,ProductNode_Float1265Output_1623);

SumNode_Float358: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float118Output_145,ProductNode_Float111Output_136,SumNode_Float358Output_1624);

ProductNode_Float1266: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v13,SumNode_Float27Output_146,ProductNode_Float1266Output_1625);

ProductNode_Float1267: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1267weight,ProductNode_Float119Output_147,ProductNode_Float1267Output_1626);

ProductNode_Float1268: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1268weight,v11,ProductNode_Float1268Output_1627);

ProductNode_Float1269: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1269weight,vb11,ProductNode_Float1269Output_1628);

SumNode_Float359: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float122Output_150,ProductNode_Float121Output_149,SumNode_Float359Output_1629);

ProductNode_Float1270: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v12,SumNode_Float28Output_151,ProductNode_Float1270Output_1630);

ProductNode_Float1271: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1271weight,ProductNode_Float123Output_152,ProductNode_Float1271Output_1631);

ProductNode_Float1272: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1272weight,v2,ProductNode_Float1272Output_1632);

ProductNode_Float1273: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1273weight,vb2,ProductNode_Float1273Output_1633);

SumNode_Float360: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float126Output_155,ProductNode_Float125Output_154,SumNode_Float360Output_1634);

ProductNode_Float1274: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float29Output_156,ProductNode_Float124Output_153,ProductNode_Float1274Output_1635);

ProductNode_Float1275: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1275weight,v11,ProductNode_Float1275Output_1636);

ProductNode_Float1276: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1276weight,vb11,ProductNode_Float1276Output_1637);

SumNode_Float361: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float129Output_159,ProductNode_Float128Output_158,SumNode_Float361Output_1638);

ProductNode_Float1277: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb12,SumNode_Float30Output_160,ProductNode_Float1277Output_1639);

ProductNode_Float1278: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1278weight,ProductNode_Float130Output_161,ProductNode_Float1278Output_1640);

ProductNode_Float1279: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1279weight,v2,ProductNode_Float1279Output_1641);

ProductNode_Float1280: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1280weight,vb2,ProductNode_Float1280Output_1642);

SumNode_Float362: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float133Output_164,ProductNode_Float132Output_163,SumNode_Float362Output_1643);

ProductNode_Float1281: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float31Output_165,ProductNode_Float131Output_162,ProductNode_Float1281Output_1644);

SumNode_Float363: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float134Output_166,ProductNode_Float127Output_157,SumNode_Float363Output_1645);

ProductNode_Float1282: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb13,SumNode_Float32Output_167,ProductNode_Float1282Output_1646);

ProductNode_Float1283: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1283weight,ProductNode_Float135Output_168,ProductNode_Float1283Output_1647);

SumNode_Float364: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float136Output_169,ProductNode_Float120Output_148,SumNode_Float364Output_1648);

ProductNode_Float1284: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v10,SumNode_Float33Output_170,ProductNode_Float1284Output_1649);

ProductNode_Float1285: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1285weight,v1,ProductNode_Float1285Output_1650);

ProductNode_Float1286: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1286weight,vb1,ProductNode_Float1286Output_1651);

SumNode_Float365: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1286Output_1651,ProductNode_Float1285Output_1650,SumNode_Float365Output_1652);

ProductNode_Float1287: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v9,SumNode_Float365Output_1652,ProductNode_Float1287Output_1653);

ProductNode_Float1288: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1288weight,ProductNode_Float1287Output_1653,ProductNode_Float1288Output_1654);

ProductNode_Float1289: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1289weight,ProductNode_Float1288Output_1654,ProductNode_Float1289Output_1655);

ProductNode_Float1290: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1290weight,v1,ProductNode_Float1290Output_1656);

ProductNode_Float1291: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1291weight,vb1,ProductNode_Float1291Output_1657);

SumNode_Float366: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1291Output_1657,ProductNode_Float1290Output_1656,SumNode_Float366Output_1658);

ProductNode_Float1292: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb9,SumNode_Float366Output_1658,ProductNode_Float1292Output_1659);

ProductNode_Float1293: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1293weight,ProductNode_Float1292Output_1659,ProductNode_Float1293Output_1660);

ProductNode_Float1294: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1294weight,ProductNode_Float1293Output_1660,ProductNode_Float1294Output_1661);

SumNode_Float367: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1294Output_1661,ProductNode_Float1289Output_1655,SumNode_Float367Output_1662);

ProductNode_Float1295: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float367Output_1662,ProductNode_Float137Output_171,ProductNode_Float1295Output_1663);

ProductNode_Float1296: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1296weight,v11,ProductNode_Float1296Output_1664);

ProductNode_Float1297: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1297weight,vb11,ProductNode_Float1297Output_1665);

SumNode_Float368: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float106Output_129,ProductNode_Float105Output_128,SumNode_Float368Output_1666);

ProductNode_Float1298: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v12,SumNode_Float23Output_130,ProductNode_Float1298Output_1667);

ProductNode_Float1299: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1299weight,ProductNode_Float107Output_131,ProductNode_Float1299Output_1668);

ProductNode_Float1300: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1300weight,v2,ProductNode_Float1300Output_1669);

ProductNode_Float1301: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1301weight,vb2,ProductNode_Float1301Output_1670);

SumNode_Float369: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float110Output_134,ProductNode_Float109Output_133,SumNode_Float369Output_1671);

ProductNode_Float1302: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float24Output_135,ProductNode_Float108Output_132,ProductNode_Float1302Output_1672);

ProductNode_Float1303: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1303weight,v11,ProductNode_Float1303Output_1673);

ProductNode_Float1304: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1304weight,vb11,ProductNode_Float1304Output_1674);

SumNode_Float370: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float113Output_138,ProductNode_Float112Output_137,SumNode_Float370Output_1675);

ProductNode_Float1305: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb12,SumNode_Float25Output_139,ProductNode_Float1305Output_1676);

ProductNode_Float1306: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1306weight,ProductNode_Float114Output_140,ProductNode_Float1306Output_1677);

ProductNode_Float1307: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1307weight,v2,ProductNode_Float1307Output_1678);

ProductNode_Float1308: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1308weight,vb2,ProductNode_Float1308Output_1679);

SumNode_Float371: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float117Output_143,ProductNode_Float116Output_142,SumNode_Float371Output_1680);

ProductNode_Float1309: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float26Output_144,ProductNode_Float115Output_141,ProductNode_Float1309Output_1681);

SumNode_Float372: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float118Output_145,ProductNode_Float111Output_136,SumNode_Float372Output_1682);

ProductNode_Float1310: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v13,SumNode_Float27Output_146,ProductNode_Float1310Output_1683);

ProductNode_Float1311: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1311weight,ProductNode_Float119Output_147,ProductNode_Float1311Output_1684);

ProductNode_Float1312: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1312weight,v11,ProductNode_Float1312Output_1685);

ProductNode_Float1313: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1313weight,vb11,ProductNode_Float1313Output_1686);

SumNode_Float373: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float122Output_150,ProductNode_Float121Output_149,SumNode_Float373Output_1687);

ProductNode_Float1314: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v12,SumNode_Float28Output_151,ProductNode_Float1314Output_1688);

ProductNode_Float1315: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1315weight,ProductNode_Float123Output_152,ProductNode_Float1315Output_1689);

ProductNode_Float1316: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1316weight,v2,ProductNode_Float1316Output_1690);

ProductNode_Float1317: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1317weight,vb2,ProductNode_Float1317Output_1691);

SumNode_Float374: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float126Output_155,ProductNode_Float125Output_154,SumNode_Float374Output_1692);

ProductNode_Float1318: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float29Output_156,ProductNode_Float124Output_153,ProductNode_Float1318Output_1693);

ProductNode_Float1319: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1319weight,v11,ProductNode_Float1319Output_1694);

ProductNode_Float1320: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1320weight,vb11,ProductNode_Float1320Output_1695);

SumNode_Float375: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float129Output_159,ProductNode_Float128Output_158,SumNode_Float375Output_1696);

ProductNode_Float1321: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb12,SumNode_Float30Output_160,ProductNode_Float1321Output_1697);

ProductNode_Float1322: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1322weight,ProductNode_Float130Output_161,ProductNode_Float1322Output_1698);

ProductNode_Float1323: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1323weight,v2,ProductNode_Float1323Output_1699);

ProductNode_Float1324: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1324weight,vb2,ProductNode_Float1324Output_1700);

SumNode_Float376: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float133Output_164,ProductNode_Float132Output_163,SumNode_Float376Output_1701);

ProductNode_Float1325: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float31Output_165,ProductNode_Float131Output_162,ProductNode_Float1325Output_1702);

SumNode_Float377: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float134Output_166,ProductNode_Float127Output_157,SumNode_Float377Output_1703);

ProductNode_Float1326: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb13,SumNode_Float32Output_167,ProductNode_Float1326Output_1704);

ProductNode_Float1327: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1327weight,ProductNode_Float135Output_168,ProductNode_Float1327Output_1705);

SumNode_Float378: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float180Output_227,ProductNode_Float164Output_206,SumNode_Float378Output_1706);

ProductNode_Float1328: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb10,SumNode_Float47Output_228,ProductNode_Float1328Output_1707);

ProductNode_Float1329: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1329weight,v1,ProductNode_Float1329Output_1708);

ProductNode_Float1330: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1330weight,vb1,ProductNode_Float1330Output_1709);

SumNode_Float379: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1330Output_1709,ProductNode_Float1329Output_1708,SumNode_Float379Output_1710);

ProductNode_Float1331: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v9,SumNode_Float379Output_1710,ProductNode_Float1331Output_1711);

ProductNode_Float1332: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1332weight,ProductNode_Float1331Output_1711,ProductNode_Float1332Output_1712);

ProductNode_Float1333: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1333weight,ProductNode_Float1332Output_1712,ProductNode_Float1333Output_1713);

ProductNode_Float1334: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1334weight,v1,ProductNode_Float1334Output_1714);

ProductNode_Float1335: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1335weight,vb1,ProductNode_Float1335Output_1715);

SumNode_Float380: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1335Output_1715,ProductNode_Float1334Output_1714,SumNode_Float380Output_1716);

ProductNode_Float1336: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb9,SumNode_Float380Output_1716,ProductNode_Float1336Output_1717);

ProductNode_Float1337: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1337weight,ProductNode_Float1336Output_1717,ProductNode_Float1337Output_1718);

ProductNode_Float1338: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1338weight,ProductNode_Float1337Output_1718,ProductNode_Float1338Output_1719);

SumNode_Float381: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1338Output_1719,ProductNode_Float1333Output_1713,SumNode_Float381Output_1720);

ProductNode_Float1339: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float381Output_1720,ProductNode_Float181Output_229,ProductNode_Float1339Output_1721);

SumNode_Float382: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1339Output_1721,ProductNode_Float1295Output_1663,SumNode_Float382Output_1722);

ProductNode_Float1340: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v15,SumNode_Float382Output_1722,ProductNode_Float1340Output_1723);

ProductNode_Float1341: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1341weight,ProductNode_Float1340Output_1723,ProductNode_Float1341Output_1724);

ProductNode_Float1342: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1342weight,v11,ProductNode_Float1342Output_1725);

ProductNode_Float1343: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1343weight,vb11,ProductNode_Float1343Output_1726);

SumNode_Float383: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float106Output_129,ProductNode_Float105Output_128,SumNode_Float383Output_1727);

ProductNode_Float1344: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v12,SumNode_Float23Output_130,ProductNode_Float1344Output_1728);

ProductNode_Float1345: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1345weight,ProductNode_Float107Output_131,ProductNode_Float1345Output_1729);

ProductNode_Float1346: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1346weight,v2,ProductNode_Float1346Output_1730);

ProductNode_Float1347: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1347weight,vb2,ProductNode_Float1347Output_1731);

SumNode_Float384: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float200Output_253,ProductNode_Float199Output_252,SumNode_Float384Output_1732);

ProductNode_Float1348: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float53Output_254,ProductNode_Float108Output_132,ProductNode_Float1348Output_1733);

ProductNode_Float1349: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1349weight,v11,ProductNode_Float1349Output_1734);

ProductNode_Float1350: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1350weight,vb11,ProductNode_Float1350Output_1735);

SumNode_Float385: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float113Output_138,ProductNode_Float112Output_137,SumNode_Float385Output_1736);

ProductNode_Float1351: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb12,SumNode_Float25Output_139,ProductNode_Float1351Output_1737);

ProductNode_Float1352: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1352weight,ProductNode_Float114Output_140,ProductNode_Float1352Output_1738);

ProductNode_Float1353: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1353weight,v2,ProductNode_Float1353Output_1739);

ProductNode_Float1354: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1354weight,vb2,ProductNode_Float1354Output_1740);

SumNode_Float386: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float207Output_262,ProductNode_Float206Output_261,SumNode_Float386Output_1741);

ProductNode_Float1355: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float55Output_263,ProductNode_Float115Output_141,ProductNode_Float1355Output_1742);

SumNode_Float387: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float208Output_264,ProductNode_Float201Output_255,SumNode_Float387Output_1743);

ProductNode_Float1356: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v13,SumNode_Float56Output_265,ProductNode_Float1356Output_1744);

ProductNode_Float1357: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1357weight,ProductNode_Float209Output_266,ProductNode_Float1357Output_1745);

ProductNode_Float1358: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1358weight,v11,ProductNode_Float1358Output_1746);

ProductNode_Float1359: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1359weight,vb11,ProductNode_Float1359Output_1747);

SumNode_Float388: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float122Output_150,ProductNode_Float121Output_149,SumNode_Float388Output_1748);

ProductNode_Float1360: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v12,SumNode_Float28Output_151,ProductNode_Float1360Output_1749);

ProductNode_Float1361: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1361weight,ProductNode_Float123Output_152,ProductNode_Float1361Output_1750);

ProductNode_Float1362: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1362weight,v2,ProductNode_Float1362Output_1751);

ProductNode_Float1363: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1363weight,vb2,ProductNode_Float1363Output_1752);

SumNode_Float389: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float216Output_274,ProductNode_Float215Output_273,SumNode_Float389Output_1753);

ProductNode_Float1364: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float58Output_275,ProductNode_Float124Output_153,ProductNode_Float1364Output_1754);

ProductNode_Float1365: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1365weight,v11,ProductNode_Float1365Output_1755);

ProductNode_Float1366: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1366weight,vb11,ProductNode_Float1366Output_1756);

SumNode_Float390: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float129Output_159,ProductNode_Float128Output_158,SumNode_Float390Output_1757);

ProductNode_Float1367: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb12,SumNode_Float30Output_160,ProductNode_Float1367Output_1758);

ProductNode_Float1368: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1368weight,ProductNode_Float130Output_161,ProductNode_Float1368Output_1759);

ProductNode_Float1369: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1369weight,v2,ProductNode_Float1369Output_1760);

ProductNode_Float1370: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1370weight,vb2,ProductNode_Float1370Output_1761);

SumNode_Float391: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float223Output_283,ProductNode_Float222Output_282,SumNode_Float391Output_1762);

ProductNode_Float1371: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float60Output_284,ProductNode_Float131Output_162,ProductNode_Float1371Output_1763);

SumNode_Float392: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float224Output_285,ProductNode_Float217Output_276,SumNode_Float392Output_1764);

ProductNode_Float1372: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb13,SumNode_Float61Output_286,ProductNode_Float1372Output_1765);

ProductNode_Float1373: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1373weight,ProductNode_Float225Output_287,ProductNode_Float1373Output_1766);

SumNode_Float393: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float226Output_288,ProductNode_Float210Output_267,SumNode_Float393Output_1767);

ProductNode_Float1374: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v10,SumNode_Float62Output_289,ProductNode_Float1374Output_1768);

ProductNode_Float1375: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1375weight,v1,ProductNode_Float1375Output_1769);

ProductNode_Float1376: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1376weight,vb1,ProductNode_Float1376Output_1770);

SumNode_Float394: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1286Output_1651,ProductNode_Float1285Output_1650,SumNode_Float394Output_1771);

ProductNode_Float1377: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v9,SumNode_Float365Output_1652,ProductNode_Float1377Output_1772);

ProductNode_Float1378: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1378weight,ProductNode_Float1287Output_1653,ProductNode_Float1378Output_1773);

ProductNode_Float1379: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1379weight,ProductNode_Float1378Output_1773,ProductNode_Float1379Output_1774);

ProductNode_Float1380: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1380weight,v1,ProductNode_Float1380Output_1775);

ProductNode_Float1381: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1381weight,vb1,ProductNode_Float1381Output_1776);

SumNode_Float395: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1291Output_1657,ProductNode_Float1290Output_1656,SumNode_Float395Output_1777);

ProductNode_Float1382: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb9,SumNode_Float366Output_1658,ProductNode_Float1382Output_1778);

ProductNode_Float1383: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1383weight,ProductNode_Float1292Output_1659,ProductNode_Float1383Output_1779);

ProductNode_Float1384: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1384weight,ProductNode_Float1383Output_1779,ProductNode_Float1384Output_1780);

SumNode_Float396: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1384Output_1780,ProductNode_Float1379Output_1774,SumNode_Float396Output_1781);

ProductNode_Float1385: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float396Output_1781,ProductNode_Float227Output_290,ProductNode_Float1385Output_1782);

ProductNode_Float1386: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1386weight,v11,ProductNode_Float1386Output_1783);

ProductNode_Float1387: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1387weight,vb11,ProductNode_Float1387Output_1784);

SumNode_Float397: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float106Output_129,ProductNode_Float105Output_128,SumNode_Float397Output_1785);

ProductNode_Float1388: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v12,SumNode_Float23Output_130,ProductNode_Float1388Output_1786);

ProductNode_Float1389: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1389weight,ProductNode_Float107Output_131,ProductNode_Float1389Output_1787);

ProductNode_Float1390: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1390weight,v2,ProductNode_Float1390Output_1788);

ProductNode_Float1391: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1391weight,vb2,ProductNode_Float1391Output_1789);

SumNode_Float398: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float200Output_253,ProductNode_Float199Output_252,SumNode_Float398Output_1790);

ProductNode_Float1392: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float53Output_254,ProductNode_Float108Output_132,ProductNode_Float1392Output_1791);

ProductNode_Float1393: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1393weight,v11,ProductNode_Float1393Output_1792);

ProductNode_Float1394: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1394weight,vb11,ProductNode_Float1394Output_1793);

SumNode_Float399: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float113Output_138,ProductNode_Float112Output_137,SumNode_Float399Output_1794);

ProductNode_Float1395: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb12,SumNode_Float25Output_139,ProductNode_Float1395Output_1795);

ProductNode_Float1396: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1396weight,ProductNode_Float114Output_140,ProductNode_Float1396Output_1796);

ProductNode_Float1397: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1397weight,v2,ProductNode_Float1397Output_1797);

ProductNode_Float1398: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1398weight,vb2,ProductNode_Float1398Output_1798);

SumNode_Float400: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float207Output_262,ProductNode_Float206Output_261,SumNode_Float400Output_1799);

ProductNode_Float1399: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float55Output_263,ProductNode_Float115Output_141,ProductNode_Float1399Output_1800);

SumNode_Float401: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float208Output_264,ProductNode_Float201Output_255,SumNode_Float401Output_1801);

ProductNode_Float1400: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v13,SumNode_Float56Output_265,ProductNode_Float1400Output_1802);

ProductNode_Float1401: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1401weight,ProductNode_Float209Output_266,ProductNode_Float1401Output_1803);

ProductNode_Float1402: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1402weight,v11,ProductNode_Float1402Output_1804);

ProductNode_Float1403: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1403weight,vb11,ProductNode_Float1403Output_1805);

SumNode_Float402: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float122Output_150,ProductNode_Float121Output_149,SumNode_Float402Output_1806);

ProductNode_Float1404: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v12,SumNode_Float28Output_151,ProductNode_Float1404Output_1807);

ProductNode_Float1405: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1405weight,ProductNode_Float123Output_152,ProductNode_Float1405Output_1808);

ProductNode_Float1406: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1406weight,v2,ProductNode_Float1406Output_1809);

ProductNode_Float1407: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1407weight,vb2,ProductNode_Float1407Output_1810);

SumNode_Float403: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float216Output_274,ProductNode_Float215Output_273,SumNode_Float403Output_1811);

ProductNode_Float1408: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float58Output_275,ProductNode_Float124Output_153,ProductNode_Float1408Output_1812);

ProductNode_Float1409: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1409weight,v11,ProductNode_Float1409Output_1813);

ProductNode_Float1410: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1410weight,vb11,ProductNode_Float1410Output_1814);

SumNode_Float404: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float129Output_159,ProductNode_Float128Output_158,SumNode_Float404Output_1815);

ProductNode_Float1411: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb12,SumNode_Float30Output_160,ProductNode_Float1411Output_1816);

ProductNode_Float1412: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1412weight,ProductNode_Float130Output_161,ProductNode_Float1412Output_1817);

ProductNode_Float1413: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1413weight,v2,ProductNode_Float1413Output_1818);

ProductNode_Float1414: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1414weight,vb2,ProductNode_Float1414Output_1819);

SumNode_Float405: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float223Output_283,ProductNode_Float222Output_282,SumNode_Float405Output_1820);

ProductNode_Float1415: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float60Output_284,ProductNode_Float131Output_162,ProductNode_Float1415Output_1821);

SumNode_Float406: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float224Output_285,ProductNode_Float217Output_276,SumNode_Float406Output_1822);

ProductNode_Float1416: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb13,SumNode_Float61Output_286,ProductNode_Float1416Output_1823);

ProductNode_Float1417: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1417weight,ProductNode_Float225Output_287,ProductNode_Float1417Output_1824);

SumNode_Float407: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float270Output_346,ProductNode_Float254Output_325,SumNode_Float407Output_1825);

ProductNode_Float1418: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb10,SumNode_Float76Output_347,ProductNode_Float1418Output_1826);

ProductNode_Float1419: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1419weight,v1,ProductNode_Float1419Output_1827);

ProductNode_Float1420: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1420weight,vb1,ProductNode_Float1420Output_1828);

SumNode_Float408: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1330Output_1709,ProductNode_Float1329Output_1708,SumNode_Float408Output_1829);

ProductNode_Float1421: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v9,SumNode_Float379Output_1710,ProductNode_Float1421Output_1830);

ProductNode_Float1422: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1422weight,ProductNode_Float1331Output_1711,ProductNode_Float1422Output_1831);

ProductNode_Float1423: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1423weight,ProductNode_Float1422Output_1831,ProductNode_Float1423Output_1832);

ProductNode_Float1424: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1424weight,v1,ProductNode_Float1424Output_1833);

ProductNode_Float1425: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1425weight,vb1,ProductNode_Float1425Output_1834);

SumNode_Float409: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1335Output_1715,ProductNode_Float1334Output_1714,SumNode_Float409Output_1835);

ProductNode_Float1426: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb9,SumNode_Float380Output_1716,ProductNode_Float1426Output_1836);

ProductNode_Float1427: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1427weight,ProductNode_Float1336Output_1717,ProductNode_Float1427Output_1837);

ProductNode_Float1428: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1428weight,ProductNode_Float1427Output_1837,ProductNode_Float1428Output_1838);

SumNode_Float410: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1428Output_1838,ProductNode_Float1423Output_1832,SumNode_Float410Output_1839);

ProductNode_Float1429: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float410Output_1839,ProductNode_Float271Output_348,ProductNode_Float1429Output_1840);

SumNode_Float411: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1429Output_1840,ProductNode_Float1385Output_1782,SumNode_Float411Output_1841);

ProductNode_Float1430: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb15,SumNode_Float411Output_1841,ProductNode_Float1430Output_1842);

ProductNode_Float1431: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1431weight,ProductNode_Float1430Output_1842,ProductNode_Float1431Output_1843);

SumNode_Float412: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1431Output_1843,ProductNode_Float1341Output_1724,SumNode_Float412Output_1844);

ProductNode_Float1432: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float412Output_1844,ProductNode_Float1251Output_1605,ProductNode_Float1432Output_1845);

ProductNode_Float1433: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1433weight,v4,ProductNode_Float1433Output_1846);

ProductNode_Float1434: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1434weight,v8,ProductNode_Float1434Output_1847);

ProductNode_Float1435: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1435weight,vb8,ProductNode_Float1435Output_1848);

SumNode_Float413: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2Output_2,ProductNode_Float1Output_1,SumNode_Float413Output_1849);

ProductNode_Float1436: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v7,SumNode_Float0Output_3,ProductNode_Float1436Output_1850);

ProductNode_Float1437: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1437weight,v3,ProductNode_Float1437Output_1851);

ProductNode_Float1438: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1438weight,ProductNode_Float4Output_5,ProductNode_Float1438Output_1852);

ProductNode_Float1439: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1439weight,ProductNode_Float5Output_6,ProductNode_Float1439Output_1853);

ProductNode_Float1440: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1440weight,vb3,ProductNode_Float1440Output_1854);

ProductNode_Float1441: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1441weight,ProductNode_Float7Output_8,ProductNode_Float1441Output_1855);

ProductNode_Float1442: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1442weight,ProductNode_Float8Output_9,ProductNode_Float1442Output_1856);

SumNode_Float414: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float9Output_10,ProductNode_Float6Output_7,SumNode_Float414Output_1857);

ProductNode_Float1443: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float1Output_11,ProductNode_Float3Output_4,ProductNode_Float1443Output_1858);

ProductNode_Float1444: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1444weight,ProductNode_Float10Output_12,ProductNode_Float1444Output_1859);

ProductNode_Float1445: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1445weight,v8,ProductNode_Float1445Output_1860);

ProductNode_Float1446: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1446weight,vb8,ProductNode_Float1446Output_1861);

SumNode_Float415: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float13Output_15,ProductNode_Float12Output_14,SumNode_Float415Output_1862);

ProductNode_Float1447: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb7,SumNode_Float2Output_16,ProductNode_Float1447Output_1863);

ProductNode_Float1448: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1448weight,v3,ProductNode_Float1448Output_1864);

ProductNode_Float1449: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1449weight,ProductNode_Float4Output_5,ProductNode_Float1449Output_1865);

ProductNode_Float1450: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1450weight,ProductNode_Float16Output_19,ProductNode_Float1450Output_1866);

ProductNode_Float1451: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1451weight,vb3,ProductNode_Float1451Output_1867);

ProductNode_Float1452: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1452weight,ProductNode_Float7Output_8,ProductNode_Float1452Output_1868);

ProductNode_Float1453: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1453weight,ProductNode_Float19Output_22,ProductNode_Float1453Output_1869);

SumNode_Float416: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float20Output_23,ProductNode_Float17Output_20,SumNode_Float416Output_1870);

ProductNode_Float1454: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float3Output_24,ProductNode_Float14Output_17,ProductNode_Float1454Output_1871);

ProductNode_Float1455: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1455weight,ProductNode_Float21Output_25,ProductNode_Float1455Output_1872);

SumNode_Float417: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float22Output_26,ProductNode_Float11Output_13,SumNode_Float417Output_1873);

ProductNode_Float1456: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float4Output_27,ProductNode_Float0Output_0,ProductNode_Float1456Output_1874);

ProductNode_Float1457: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1457weight,ProductNode_Float23Output_28,ProductNode_Float1457Output_1875);

ProductNode_Float1458: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1458weight,vb4,ProductNode_Float1458Output_1876);

ProductNode_Float1459: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1459weight,v8,ProductNode_Float1459Output_1877);

ProductNode_Float1460: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1460weight,vb8,ProductNode_Float1460Output_1878);

SumNode_Float418: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float27Output_32,ProductNode_Float26Output_31,SumNode_Float418Output_1879);

ProductNode_Float1461: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v7,SumNode_Float5Output_33,ProductNode_Float1461Output_1880);

ProductNode_Float1462: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1462weight,v3,ProductNode_Float1462Output_1881);

ProductNode_Float1463: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1463weight,ProductNode_Float29Output_35,ProductNode_Float1463Output_1882);

ProductNode_Float1464: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1464weight,ProductNode_Float30Output_36,ProductNode_Float1464Output_1883);

ProductNode_Float1465: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1465weight,vb3,ProductNode_Float1465Output_1884);

ProductNode_Float1466: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1466weight,ProductNode_Float32Output_38,ProductNode_Float1466Output_1885);

ProductNode_Float1467: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1467weight,ProductNode_Float33Output_39,ProductNode_Float1467Output_1886);

SumNode_Float419: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float34Output_40,ProductNode_Float31Output_37,SumNode_Float419Output_1887);

ProductNode_Float1468: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float6Output_41,ProductNode_Float28Output_34,ProductNode_Float1468Output_1888);

ProductNode_Float1469: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1469weight,ProductNode_Float35Output_42,ProductNode_Float1469Output_1889);

ProductNode_Float1470: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1470weight,v8,ProductNode_Float1470Output_1890);

ProductNode_Float1471: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1471weight,vb8,ProductNode_Float1471Output_1891);

SumNode_Float420: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float38Output_45,ProductNode_Float37Output_44,SumNode_Float420Output_1892);

ProductNode_Float1472: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb7,SumNode_Float7Output_46,ProductNode_Float1472Output_1893);

ProductNode_Float1473: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1473weight,v3,ProductNode_Float1473Output_1894);

ProductNode_Float1474: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1474weight,ProductNode_Float29Output_35,ProductNode_Float1474Output_1895);

ProductNode_Float1475: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1475weight,ProductNode_Float41Output_49,ProductNode_Float1475Output_1896);

ProductNode_Float1476: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1476weight,vb3,ProductNode_Float1476Output_1897);

ProductNode_Float1477: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1477weight,ProductNode_Float32Output_38,ProductNode_Float1477Output_1898);

ProductNode_Float1478: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1478weight,ProductNode_Float44Output_52,ProductNode_Float1478Output_1899);

SumNode_Float421: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float45Output_53,ProductNode_Float42Output_50,SumNode_Float421Output_1900);

ProductNode_Float1479: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float8Output_54,ProductNode_Float39Output_47,ProductNode_Float1479Output_1901);

ProductNode_Float1480: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1480weight,ProductNode_Float46Output_55,ProductNode_Float1480Output_1902);

SumNode_Float422: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float47Output_56,ProductNode_Float36Output_43,SumNode_Float422Output_1903);

ProductNode_Float1481: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float9Output_57,ProductNode_Float25Output_30,ProductNode_Float1481Output_1904);

ProductNode_Float1482: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1482weight,ProductNode_Float48Output_58,ProductNode_Float1482Output_1905);

SumNode_Float423: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float335Output_427,ProductNode_Float310Output_397,SumNode_Float423Output_1906);

ProductNode_Float1483: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v5,SumNode_Float92Output_428,ProductNode_Float1483Output_1907);

ProductNode_Float1484: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1484weight,ProductNode_Float336Output_429,ProductNode_Float1484Output_1908);

ProductNode_Float1485: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1485weight,v4,ProductNode_Float1485Output_1909);

ProductNode_Float1486: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1486weight,v8,ProductNode_Float1486Output_1910);

ProductNode_Float1487: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1487weight,vb8,ProductNode_Float1487Output_1911);

SumNode_Float424: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float54Output_65,ProductNode_Float53Output_64,SumNode_Float424Output_1912);

ProductNode_Float1488: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v7,SumNode_Float11Output_66,ProductNode_Float1488Output_1913);

ProductNode_Float1489: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1489weight,v3,ProductNode_Float1489Output_1914);

ProductNode_Float1490: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1490weight,ProductNode_Float4Output_5,ProductNode_Float1490Output_1915);

ProductNode_Float1491: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1491weight,ProductNode_Float5Output_6,ProductNode_Float1491Output_1916);

ProductNode_Float1492: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1492weight,vb3,ProductNode_Float1492Output_1917);

ProductNode_Float1493: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1493weight,ProductNode_Float7Output_8,ProductNode_Float1493Output_1918);

ProductNode_Float1494: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1494weight,ProductNode_Float8Output_9,ProductNode_Float1494Output_1919);

SumNode_Float425: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float61Output_73,ProductNode_Float58Output_70,SumNode_Float425Output_1920);

ProductNode_Float1495: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float12Output_74,ProductNode_Float55Output_67,ProductNode_Float1495Output_1921);

ProductNode_Float1496: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1496weight,ProductNode_Float62Output_75,ProductNode_Float1496Output_1922);

ProductNode_Float1497: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1497weight,v8,ProductNode_Float1497Output_1923);

ProductNode_Float1498: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1498weight,vb8,ProductNode_Float1498Output_1924);

SumNode_Float426: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float65Output_78,ProductNode_Float64Output_77,SumNode_Float426Output_1925);

ProductNode_Float1499: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb7,SumNode_Float13Output_79,ProductNode_Float1499Output_1926);

ProductNode_Float1500: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1500weight,v3,ProductNode_Float1500Output_1927);

ProductNode_Float1501: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1501weight,ProductNode_Float4Output_5,ProductNode_Float1501Output_1928);

ProductNode_Float1502: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1502weight,ProductNode_Float16Output_19,ProductNode_Float1502Output_1929);

ProductNode_Float1503: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1503weight,vb3,ProductNode_Float1503Output_1930);

ProductNode_Float1504: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1504weight,ProductNode_Float7Output_8,ProductNode_Float1504Output_1931);

ProductNode_Float1505: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1505weight,ProductNode_Float19Output_22,ProductNode_Float1505Output_1932);

SumNode_Float427: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float72Output_86,ProductNode_Float69Output_83,SumNode_Float427Output_1933);

ProductNode_Float1506: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float14Output_87,ProductNode_Float66Output_80,ProductNode_Float1506Output_1934);

ProductNode_Float1507: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1507weight,ProductNode_Float73Output_88,ProductNode_Float1507Output_1935);

SumNode_Float428: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float74Output_89,ProductNode_Float63Output_76,SumNode_Float428Output_1936);

ProductNode_Float1508: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float15Output_90,ProductNode_Float0Output_0,ProductNode_Float1508Output_1937);

ProductNode_Float1509: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1509weight,ProductNode_Float75Output_91,ProductNode_Float1509Output_1938);

ProductNode_Float1510: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1510weight,vb4,ProductNode_Float1510Output_1939);

ProductNode_Float1511: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1511weight,v8,ProductNode_Float1511Output_1940);

ProductNode_Float1512: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1512weight,vb8,ProductNode_Float1512Output_1941);

SumNode_Float429: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float79Output_95,ProductNode_Float78Output_94,SumNode_Float429Output_1942);

ProductNode_Float1513: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v7,SumNode_Float16Output_96,ProductNode_Float1513Output_1943);

ProductNode_Float1514: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1514weight,v3,ProductNode_Float1514Output_1944);

ProductNode_Float1515: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1515weight,ProductNode_Float29Output_35,ProductNode_Float1515Output_1945);

ProductNode_Float1516: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1516weight,ProductNode_Float30Output_36,ProductNode_Float1516Output_1946);

ProductNode_Float1517: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1517weight,vb3,ProductNode_Float1517Output_1947);

ProductNode_Float1518: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1518weight,ProductNode_Float32Output_38,ProductNode_Float1518Output_1948);

ProductNode_Float1519: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1519weight,ProductNode_Float33Output_39,ProductNode_Float1519Output_1949);

SumNode_Float430: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float86Output_103,ProductNode_Float83Output_100,SumNode_Float430Output_1950);

ProductNode_Float1520: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float17Output_104,ProductNode_Float80Output_97,ProductNode_Float1520Output_1951);

ProductNode_Float1521: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1521weight,ProductNode_Float87Output_105,ProductNode_Float1521Output_1952);

ProductNode_Float1522: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1522weight,v8,ProductNode_Float1522Output_1953);

ProductNode_Float1523: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1523weight,vb8,ProductNode_Float1523Output_1954);

SumNode_Float431: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float90Output_108,ProductNode_Float89Output_107,SumNode_Float431Output_1955);

ProductNode_Float1524: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb7,SumNode_Float18Output_109,ProductNode_Float1524Output_1956);

ProductNode_Float1525: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1525weight,v3,ProductNode_Float1525Output_1957);

ProductNode_Float1526: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1526weight,ProductNode_Float29Output_35,ProductNode_Float1526Output_1958);

ProductNode_Float1527: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1527weight,ProductNode_Float41Output_49,ProductNode_Float1527Output_1959);

ProductNode_Float1528: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1528weight,vb3,ProductNode_Float1528Output_1960);

ProductNode_Float1529: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1529weight,ProductNode_Float32Output_38,ProductNode_Float1529Output_1961);

ProductNode_Float1530: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1530weight,ProductNode_Float44Output_52,ProductNode_Float1530Output_1962);

SumNode_Float432: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float97Output_116,ProductNode_Float94Output_113,SumNode_Float432Output_1963);

ProductNode_Float1531: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float19Output_117,ProductNode_Float91Output_110,ProductNode_Float1531Output_1964);

ProductNode_Float1532: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1532weight,ProductNode_Float98Output_118,ProductNode_Float1532Output_1965);

SumNode_Float433: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float99Output_119,ProductNode_Float88Output_106,SumNode_Float433Output_1966);

ProductNode_Float1533: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float20Output_120,ProductNode_Float25Output_30,ProductNode_Float1533Output_1967);

ProductNode_Float1534: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1534weight,ProductNode_Float100Output_121,ProductNode_Float1534Output_1968);

SumNode_Float434: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float387Output_490,ProductNode_Float362Output_460,SumNode_Float434Output_1969);

ProductNode_Float1535: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb5,SumNode_Float103Output_491,ProductNode_Float1535Output_1970);

ProductNode_Float1536: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1536weight,ProductNode_Float388Output_492,ProductNode_Float1536Output_1971);

SumNode_Float435: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1536Output_1971,ProductNode_Float1484Output_1908,SumNode_Float435Output_1972);

ProductNode_Float1537: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb16,SumNode_Float435Output_1972,ProductNode_Float1537Output_1973);

ProductNode_Float1538: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1538weight,v11,ProductNode_Float1538Output_1974);

ProductNode_Float1539: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1539weight,vb11,ProductNode_Float1539Output_1975);

SumNode_Float436: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float106Output_129,ProductNode_Float105Output_128,SumNode_Float436Output_1976);

ProductNode_Float1540: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v12,SumNode_Float23Output_130,ProductNode_Float1540Output_1977);

ProductNode_Float1541: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1541weight,ProductNode_Float107Output_131,ProductNode_Float1541Output_1978);

ProductNode_Float1542: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1542weight,v2,ProductNode_Float1542Output_1979);

ProductNode_Float1543: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1543weight,vb2,ProductNode_Float1543Output_1980);

SumNode_Float437: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float110Output_134,ProductNode_Float109Output_133,SumNode_Float437Output_1981);

ProductNode_Float1544: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float24Output_135,ProductNode_Float108Output_132,ProductNode_Float1544Output_1982);

ProductNode_Float1545: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1545weight,v11,ProductNode_Float1545Output_1983);

ProductNode_Float1546: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1546weight,vb11,ProductNode_Float1546Output_1984);

SumNode_Float438: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float113Output_138,ProductNode_Float112Output_137,SumNode_Float438Output_1985);

ProductNode_Float1547: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb12,SumNode_Float25Output_139,ProductNode_Float1547Output_1986);

ProductNode_Float1548: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1548weight,ProductNode_Float114Output_140,ProductNode_Float1548Output_1987);

ProductNode_Float1549: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1549weight,v2,ProductNode_Float1549Output_1988);

ProductNode_Float1550: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1550weight,vb2,ProductNode_Float1550Output_1989);

SumNode_Float439: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float117Output_143,ProductNode_Float116Output_142,SumNode_Float439Output_1990);

ProductNode_Float1551: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float26Output_144,ProductNode_Float115Output_141,ProductNode_Float1551Output_1991);

SumNode_Float440: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float118Output_145,ProductNode_Float111Output_136,SumNode_Float440Output_1992);

ProductNode_Float1552: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v13,SumNode_Float27Output_146,ProductNode_Float1552Output_1993);

ProductNode_Float1553: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1553weight,ProductNode_Float119Output_147,ProductNode_Float1553Output_1994);

ProductNode_Float1554: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1554weight,v11,ProductNode_Float1554Output_1995);

ProductNode_Float1555: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1555weight,vb11,ProductNode_Float1555Output_1996);

SumNode_Float441: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float122Output_150,ProductNode_Float121Output_149,SumNode_Float441Output_1997);

ProductNode_Float1556: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v12,SumNode_Float28Output_151,ProductNode_Float1556Output_1998);

ProductNode_Float1557: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1557weight,ProductNode_Float123Output_152,ProductNode_Float1557Output_1999);

ProductNode_Float1558: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1558weight,v2,ProductNode_Float1558Output_2000);

ProductNode_Float1559: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1559weight,vb2,ProductNode_Float1559Output_2001);

SumNode_Float442: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float126Output_155,ProductNode_Float125Output_154,SumNode_Float442Output_2002);

ProductNode_Float1560: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float29Output_156,ProductNode_Float124Output_153,ProductNode_Float1560Output_2003);

ProductNode_Float1561: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1561weight,v11,ProductNode_Float1561Output_2004);

ProductNode_Float1562: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1562weight,vb11,ProductNode_Float1562Output_2005);

SumNode_Float443: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float129Output_159,ProductNode_Float128Output_158,SumNode_Float443Output_2006);

ProductNode_Float1563: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb12,SumNode_Float30Output_160,ProductNode_Float1563Output_2007);

ProductNode_Float1564: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1564weight,ProductNode_Float130Output_161,ProductNode_Float1564Output_2008);

ProductNode_Float1565: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1565weight,v2,ProductNode_Float1565Output_2009);

ProductNode_Float1566: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1566weight,vb2,ProductNode_Float1566Output_2010);

SumNode_Float444: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float133Output_164,ProductNode_Float132Output_163,SumNode_Float444Output_2011);

ProductNode_Float1567: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float31Output_165,ProductNode_Float131Output_162,ProductNode_Float1567Output_2012);

SumNode_Float445: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float134Output_166,ProductNode_Float127Output_157,SumNode_Float445Output_2013);

ProductNode_Float1568: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb13,SumNode_Float32Output_167,ProductNode_Float1568Output_2014);

ProductNode_Float1569: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1569weight,ProductNode_Float135Output_168,ProductNode_Float1569Output_2015);

SumNode_Float446: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float136Output_169,ProductNode_Float120Output_148,SumNode_Float446Output_2016);

ProductNode_Float1570: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v10,SumNode_Float33Output_170,ProductNode_Float1570Output_2017);

ProductNode_Float1571: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1571weight,v1,ProductNode_Float1571Output_2018);

ProductNode_Float1572: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1572weight,vb1,ProductNode_Float1572Output_2019);

SumNode_Float447: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1286Output_1651,ProductNode_Float1285Output_1650,SumNode_Float447Output_2020);

ProductNode_Float1573: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v9,SumNode_Float365Output_1652,ProductNode_Float1573Output_2021);

ProductNode_Float1574: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1574weight,ProductNode_Float1287Output_1653,ProductNode_Float1574Output_2022);

ProductNode_Float1575: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1575weight,ProductNode_Float1288Output_1654,ProductNode_Float1575Output_2023);

ProductNode_Float1576: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1576weight,v1,ProductNode_Float1576Output_2024);

ProductNode_Float1577: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1577weight,vb1,ProductNode_Float1577Output_2025);

SumNode_Float448: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1291Output_1657,ProductNode_Float1290Output_1656,SumNode_Float448Output_2026);

ProductNode_Float1578: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb9,SumNode_Float366Output_1658,ProductNode_Float1578Output_2027);

ProductNode_Float1579: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1579weight,ProductNode_Float1292Output_1659,ProductNode_Float1579Output_2028);

ProductNode_Float1580: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1580weight,ProductNode_Float1293Output_1660,ProductNode_Float1580Output_2029);

SumNode_Float449: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1294Output_1661,ProductNode_Float1289Output_1655,SumNode_Float449Output_2030);

ProductNode_Float1581: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float367Output_1662,ProductNode_Float137Output_171,ProductNode_Float1581Output_2031);

ProductNode_Float1582: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1582weight,v11,ProductNode_Float1582Output_2032);

ProductNode_Float1583: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1583weight,vb11,ProductNode_Float1583Output_2033);

SumNode_Float450: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float106Output_129,ProductNode_Float105Output_128,SumNode_Float450Output_2034);

ProductNode_Float1584: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v12,SumNode_Float23Output_130,ProductNode_Float1584Output_2035);

ProductNode_Float1585: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1585weight,ProductNode_Float107Output_131,ProductNode_Float1585Output_2036);

ProductNode_Float1586: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1586weight,v2,ProductNode_Float1586Output_2037);

ProductNode_Float1587: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1587weight,vb2,ProductNode_Float1587Output_2038);

SumNode_Float451: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float110Output_134,ProductNode_Float109Output_133,SumNode_Float451Output_2039);

ProductNode_Float1588: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float24Output_135,ProductNode_Float108Output_132,ProductNode_Float1588Output_2040);

ProductNode_Float1589: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1589weight,v11,ProductNode_Float1589Output_2041);

ProductNode_Float1590: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1590weight,vb11,ProductNode_Float1590Output_2042);

SumNode_Float452: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float113Output_138,ProductNode_Float112Output_137,SumNode_Float452Output_2043);

ProductNode_Float1591: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb12,SumNode_Float25Output_139,ProductNode_Float1591Output_2044);

ProductNode_Float1592: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1592weight,ProductNode_Float114Output_140,ProductNode_Float1592Output_2045);

ProductNode_Float1593: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1593weight,v2,ProductNode_Float1593Output_2046);

ProductNode_Float1594: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1594weight,vb2,ProductNode_Float1594Output_2047);

SumNode_Float453: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float117Output_143,ProductNode_Float116Output_142,SumNode_Float453Output_2048);

ProductNode_Float1595: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float26Output_144,ProductNode_Float115Output_141,ProductNode_Float1595Output_2049);

SumNode_Float454: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float118Output_145,ProductNode_Float111Output_136,SumNode_Float454Output_2050);

ProductNode_Float1596: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v13,SumNode_Float27Output_146,ProductNode_Float1596Output_2051);

ProductNode_Float1597: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1597weight,ProductNode_Float119Output_147,ProductNode_Float1597Output_2052);

ProductNode_Float1598: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1598weight,v11,ProductNode_Float1598Output_2053);

ProductNode_Float1599: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1599weight,vb11,ProductNode_Float1599Output_2054);

SumNode_Float455: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float122Output_150,ProductNode_Float121Output_149,SumNode_Float455Output_2055);

ProductNode_Float1600: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v12,SumNode_Float28Output_151,ProductNode_Float1600Output_2056);

ProductNode_Float1601: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1601weight,ProductNode_Float123Output_152,ProductNode_Float1601Output_2057);

ProductNode_Float1602: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1602weight,v2,ProductNode_Float1602Output_2058);

ProductNode_Float1603: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1603weight,vb2,ProductNode_Float1603Output_2059);

SumNode_Float456: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float126Output_155,ProductNode_Float125Output_154,SumNode_Float456Output_2060);

ProductNode_Float1604: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float29Output_156,ProductNode_Float124Output_153,ProductNode_Float1604Output_2061);

ProductNode_Float1605: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1605weight,v11,ProductNode_Float1605Output_2062);

ProductNode_Float1606: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1606weight,vb11,ProductNode_Float1606Output_2063);

SumNode_Float457: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float129Output_159,ProductNode_Float128Output_158,SumNode_Float457Output_2064);

ProductNode_Float1607: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb12,SumNode_Float30Output_160,ProductNode_Float1607Output_2065);

ProductNode_Float1608: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1608weight,ProductNode_Float130Output_161,ProductNode_Float1608Output_2066);

ProductNode_Float1609: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1609weight,v2,ProductNode_Float1609Output_2067);

ProductNode_Float1610: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1610weight,vb2,ProductNode_Float1610Output_2068);

SumNode_Float458: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float133Output_164,ProductNode_Float132Output_163,SumNode_Float458Output_2069);

ProductNode_Float1611: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float31Output_165,ProductNode_Float131Output_162,ProductNode_Float1611Output_2070);

SumNode_Float459: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float134Output_166,ProductNode_Float127Output_157,SumNode_Float459Output_2071);

ProductNode_Float1612: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb13,SumNode_Float32Output_167,ProductNode_Float1612Output_2072);

ProductNode_Float1613: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1613weight,ProductNode_Float135Output_168,ProductNode_Float1613Output_2073);

SumNode_Float460: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float180Output_227,ProductNode_Float164Output_206,SumNode_Float460Output_2074);

ProductNode_Float1614: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb10,SumNode_Float47Output_228,ProductNode_Float1614Output_2075);

ProductNode_Float1615: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1615weight,v1,ProductNode_Float1615Output_2076);

ProductNode_Float1616: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1616weight,vb1,ProductNode_Float1616Output_2077);

SumNode_Float461: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1330Output_1709,ProductNode_Float1329Output_1708,SumNode_Float461Output_2078);

ProductNode_Float1617: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v9,SumNode_Float379Output_1710,ProductNode_Float1617Output_2079);

ProductNode_Float1618: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1618weight,ProductNode_Float1331Output_1711,ProductNode_Float1618Output_2080);

ProductNode_Float1619: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1619weight,ProductNode_Float1332Output_1712,ProductNode_Float1619Output_2081);

ProductNode_Float1620: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1620weight,v1,ProductNode_Float1620Output_2082);

ProductNode_Float1621: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1621weight,vb1,ProductNode_Float1621Output_2083);

SumNode_Float462: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1335Output_1715,ProductNode_Float1334Output_1714,SumNode_Float462Output_2084);

ProductNode_Float1622: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb9,SumNode_Float380Output_1716,ProductNode_Float1622Output_2085);

ProductNode_Float1623: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1623weight,ProductNode_Float1336Output_1717,ProductNode_Float1623Output_2086);

ProductNode_Float1624: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1624weight,ProductNode_Float1337Output_1718,ProductNode_Float1624Output_2087);

SumNode_Float463: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1338Output_1719,ProductNode_Float1333Output_1713,SumNode_Float463Output_2088);

ProductNode_Float1625: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float381Output_1720,ProductNode_Float181Output_229,ProductNode_Float1625Output_2089);

SumNode_Float464: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1339Output_1721,ProductNode_Float1295Output_1663,SumNode_Float464Output_2090);

ProductNode_Float1626: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v15,SumNode_Float382Output_1722,ProductNode_Float1626Output_2091);

ProductNode_Float1627: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1627weight,ProductNode_Float1340Output_1723,ProductNode_Float1627Output_2092);

ProductNode_Float1628: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1628weight,v11,ProductNode_Float1628Output_2093);

ProductNode_Float1629: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1629weight,vb11,ProductNode_Float1629Output_2094);

SumNode_Float465: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float106Output_129,ProductNode_Float105Output_128,SumNode_Float465Output_2095);

ProductNode_Float1630: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v12,SumNode_Float23Output_130,ProductNode_Float1630Output_2096);

ProductNode_Float1631: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1631weight,ProductNode_Float107Output_131,ProductNode_Float1631Output_2097);

ProductNode_Float1632: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1632weight,v2,ProductNode_Float1632Output_2098);

ProductNode_Float1633: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1633weight,vb2,ProductNode_Float1633Output_2099);

SumNode_Float466: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float200Output_253,ProductNode_Float199Output_252,SumNode_Float466Output_2100);

ProductNode_Float1634: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float53Output_254,ProductNode_Float108Output_132,ProductNode_Float1634Output_2101);

ProductNode_Float1635: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1635weight,v11,ProductNode_Float1635Output_2102);

ProductNode_Float1636: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1636weight,vb11,ProductNode_Float1636Output_2103);

SumNode_Float467: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float113Output_138,ProductNode_Float112Output_137,SumNode_Float467Output_2104);

ProductNode_Float1637: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb12,SumNode_Float25Output_139,ProductNode_Float1637Output_2105);

ProductNode_Float1638: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1638weight,ProductNode_Float114Output_140,ProductNode_Float1638Output_2106);

ProductNode_Float1639: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1639weight,v2,ProductNode_Float1639Output_2107);

ProductNode_Float1640: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1640weight,vb2,ProductNode_Float1640Output_2108);

SumNode_Float468: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float207Output_262,ProductNode_Float206Output_261,SumNode_Float468Output_2109);

ProductNode_Float1641: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float55Output_263,ProductNode_Float115Output_141,ProductNode_Float1641Output_2110);

SumNode_Float469: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float208Output_264,ProductNode_Float201Output_255,SumNode_Float469Output_2111);

ProductNode_Float1642: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v13,SumNode_Float56Output_265,ProductNode_Float1642Output_2112);

ProductNode_Float1643: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1643weight,ProductNode_Float209Output_266,ProductNode_Float1643Output_2113);

ProductNode_Float1644: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1644weight,v11,ProductNode_Float1644Output_2114);

ProductNode_Float1645: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1645weight,vb11,ProductNode_Float1645Output_2115);

SumNode_Float470: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float122Output_150,ProductNode_Float121Output_149,SumNode_Float470Output_2116);

ProductNode_Float1646: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v12,SumNode_Float28Output_151,ProductNode_Float1646Output_2117);

ProductNode_Float1647: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1647weight,ProductNode_Float123Output_152,ProductNode_Float1647Output_2118);

ProductNode_Float1648: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1648weight,v2,ProductNode_Float1648Output_2119);

ProductNode_Float1649: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1649weight,vb2,ProductNode_Float1649Output_2120);

SumNode_Float471: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float216Output_274,ProductNode_Float215Output_273,SumNode_Float471Output_2121);

ProductNode_Float1650: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float58Output_275,ProductNode_Float124Output_153,ProductNode_Float1650Output_2122);

ProductNode_Float1651: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1651weight,v11,ProductNode_Float1651Output_2123);

ProductNode_Float1652: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1652weight,vb11,ProductNode_Float1652Output_2124);

SumNode_Float472: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float129Output_159,ProductNode_Float128Output_158,SumNode_Float472Output_2125);

ProductNode_Float1653: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb12,SumNode_Float30Output_160,ProductNode_Float1653Output_2126);

ProductNode_Float1654: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1654weight,ProductNode_Float130Output_161,ProductNode_Float1654Output_2127);

ProductNode_Float1655: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1655weight,v2,ProductNode_Float1655Output_2128);

ProductNode_Float1656: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1656weight,vb2,ProductNode_Float1656Output_2129);

SumNode_Float473: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float223Output_283,ProductNode_Float222Output_282,SumNode_Float473Output_2130);

ProductNode_Float1657: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float60Output_284,ProductNode_Float131Output_162,ProductNode_Float1657Output_2131);

SumNode_Float474: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float224Output_285,ProductNode_Float217Output_276,SumNode_Float474Output_2132);

ProductNode_Float1658: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb13,SumNode_Float61Output_286,ProductNode_Float1658Output_2133);

ProductNode_Float1659: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1659weight,ProductNode_Float225Output_287,ProductNode_Float1659Output_2134);

SumNode_Float475: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float226Output_288,ProductNode_Float210Output_267,SumNode_Float475Output_2135);

ProductNode_Float1660: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v10,SumNode_Float62Output_289,ProductNode_Float1660Output_2136);

ProductNode_Float1661: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1661weight,v1,ProductNode_Float1661Output_2137);

ProductNode_Float1662: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1662weight,vb1,ProductNode_Float1662Output_2138);

SumNode_Float476: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1286Output_1651,ProductNode_Float1285Output_1650,SumNode_Float476Output_2139);

ProductNode_Float1663: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v9,SumNode_Float365Output_1652,ProductNode_Float1663Output_2140);

ProductNode_Float1664: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1664weight,ProductNode_Float1287Output_1653,ProductNode_Float1664Output_2141);

ProductNode_Float1665: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1665weight,ProductNode_Float1378Output_1773,ProductNode_Float1665Output_2142);

ProductNode_Float1666: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1666weight,v1,ProductNode_Float1666Output_2143);

ProductNode_Float1667: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1667weight,vb1,ProductNode_Float1667Output_2144);

SumNode_Float477: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1291Output_1657,ProductNode_Float1290Output_1656,SumNode_Float477Output_2145);

ProductNode_Float1668: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb9,SumNode_Float366Output_1658,ProductNode_Float1668Output_2146);

ProductNode_Float1669: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1669weight,ProductNode_Float1292Output_1659,ProductNode_Float1669Output_2147);

ProductNode_Float1670: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1670weight,ProductNode_Float1383Output_1779,ProductNode_Float1670Output_2148);

SumNode_Float478: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1384Output_1780,ProductNode_Float1379Output_1774,SumNode_Float478Output_2149);

ProductNode_Float1671: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float396Output_1781,ProductNode_Float227Output_290,ProductNode_Float1671Output_2150);

ProductNode_Float1672: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1672weight,v11,ProductNode_Float1672Output_2151);

ProductNode_Float1673: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1673weight,vb11,ProductNode_Float1673Output_2152);

SumNode_Float479: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float106Output_129,ProductNode_Float105Output_128,SumNode_Float479Output_2153);

ProductNode_Float1674: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v12,SumNode_Float23Output_130,ProductNode_Float1674Output_2154);

ProductNode_Float1675: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1675weight,ProductNode_Float107Output_131,ProductNode_Float1675Output_2155);

ProductNode_Float1676: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1676weight,v2,ProductNode_Float1676Output_2156);

ProductNode_Float1677: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1677weight,vb2,ProductNode_Float1677Output_2157);

SumNode_Float480: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float200Output_253,ProductNode_Float199Output_252,SumNode_Float480Output_2158);

ProductNode_Float1678: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float53Output_254,ProductNode_Float108Output_132,ProductNode_Float1678Output_2159);

ProductNode_Float1679: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1679weight,v11,ProductNode_Float1679Output_2160);

ProductNode_Float1680: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1680weight,vb11,ProductNode_Float1680Output_2161);

SumNode_Float481: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float113Output_138,ProductNode_Float112Output_137,SumNode_Float481Output_2162);

ProductNode_Float1681: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb12,SumNode_Float25Output_139,ProductNode_Float1681Output_2163);

ProductNode_Float1682: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1682weight,ProductNode_Float114Output_140,ProductNode_Float1682Output_2164);

ProductNode_Float1683: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1683weight,v2,ProductNode_Float1683Output_2165);

ProductNode_Float1684: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1684weight,vb2,ProductNode_Float1684Output_2166);

SumNode_Float482: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float207Output_262,ProductNode_Float206Output_261,SumNode_Float482Output_2167);

ProductNode_Float1685: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float55Output_263,ProductNode_Float115Output_141,ProductNode_Float1685Output_2168);

SumNode_Float483: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float208Output_264,ProductNode_Float201Output_255,SumNode_Float483Output_2169);

ProductNode_Float1686: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v13,SumNode_Float56Output_265,ProductNode_Float1686Output_2170);

ProductNode_Float1687: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1687weight,ProductNode_Float209Output_266,ProductNode_Float1687Output_2171);

ProductNode_Float1688: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1688weight,v11,ProductNode_Float1688Output_2172);

ProductNode_Float1689: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1689weight,vb11,ProductNode_Float1689Output_2173);

SumNode_Float484: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float122Output_150,ProductNode_Float121Output_149,SumNode_Float484Output_2174);

ProductNode_Float1690: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v12,SumNode_Float28Output_151,ProductNode_Float1690Output_2175);

ProductNode_Float1691: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1691weight,ProductNode_Float123Output_152,ProductNode_Float1691Output_2176);

ProductNode_Float1692: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1692weight,v2,ProductNode_Float1692Output_2177);

ProductNode_Float1693: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1693weight,vb2,ProductNode_Float1693Output_2178);

SumNode_Float485: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float216Output_274,ProductNode_Float215Output_273,SumNode_Float485Output_2179);

ProductNode_Float1694: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float58Output_275,ProductNode_Float124Output_153,ProductNode_Float1694Output_2180);

ProductNode_Float1695: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1695weight,v11,ProductNode_Float1695Output_2181);

ProductNode_Float1696: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1696weight,vb11,ProductNode_Float1696Output_2182);

SumNode_Float486: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float129Output_159,ProductNode_Float128Output_158,SumNode_Float486Output_2183);

ProductNode_Float1697: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb12,SumNode_Float30Output_160,ProductNode_Float1697Output_2184);

ProductNode_Float1698: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1698weight,ProductNode_Float130Output_161,ProductNode_Float1698Output_2185);

ProductNode_Float1699: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1699weight,v2,ProductNode_Float1699Output_2186);

ProductNode_Float1700: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1700weight,vb2,ProductNode_Float1700Output_2187);

SumNode_Float487: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float223Output_283,ProductNode_Float222Output_282,SumNode_Float487Output_2188);

ProductNode_Float1701: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float60Output_284,ProductNode_Float131Output_162,ProductNode_Float1701Output_2189);

SumNode_Float488: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float224Output_285,ProductNode_Float217Output_276,SumNode_Float488Output_2190);

ProductNode_Float1702: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb13,SumNode_Float61Output_286,ProductNode_Float1702Output_2191);

ProductNode_Float1703: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1703weight,ProductNode_Float225Output_287,ProductNode_Float1703Output_2192);

SumNode_Float489: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float270Output_346,ProductNode_Float254Output_325,SumNode_Float489Output_2193);

ProductNode_Float1704: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb10,SumNode_Float76Output_347,ProductNode_Float1704Output_2194);

ProductNode_Float1705: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1705weight,v1,ProductNode_Float1705Output_2195);

ProductNode_Float1706: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1706weight,vb1,ProductNode_Float1706Output_2196);

SumNode_Float490: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1330Output_1709,ProductNode_Float1329Output_1708,SumNode_Float490Output_2197);

ProductNode_Float1707: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v9,SumNode_Float379Output_1710,ProductNode_Float1707Output_2198);

ProductNode_Float1708: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1708weight,ProductNode_Float1331Output_1711,ProductNode_Float1708Output_2199);

ProductNode_Float1709: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1709weight,ProductNode_Float1422Output_1831,ProductNode_Float1709Output_2200);

ProductNode_Float1710: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1710weight,v1,ProductNode_Float1710Output_2201);

ProductNode_Float1711: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1711weight,vb1,ProductNode_Float1711Output_2202);

SumNode_Float491: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1335Output_1715,ProductNode_Float1334Output_1714,SumNode_Float491Output_2203);

ProductNode_Float1712: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb9,SumNode_Float380Output_1716,ProductNode_Float1712Output_2204);

ProductNode_Float1713: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1713weight,ProductNode_Float1336Output_1717,ProductNode_Float1713Output_2205);

ProductNode_Float1714: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1714weight,ProductNode_Float1427Output_1837,ProductNode_Float1714Output_2206);

SumNode_Float492: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1428Output_1838,ProductNode_Float1423Output_1832,SumNode_Float492Output_2207);

ProductNode_Float1715: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float410Output_1839,ProductNode_Float271Output_348,ProductNode_Float1715Output_2208);

SumNode_Float493: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1429Output_1840,ProductNode_Float1385Output_1782,SumNode_Float493Output_2209);

ProductNode_Float1716: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb15,SumNode_Float411Output_1841,ProductNode_Float1716Output_2210);

ProductNode_Float1717: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1717weight,ProductNode_Float1430Output_1842,ProductNode_Float1717Output_2211);

SumNode_Float494: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1717Output_2211,ProductNode_Float1627Output_2092,SumNode_Float494Output_2212);

ProductNode_Float1718: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float494Output_2212,ProductNode_Float1537Output_1973,ProductNode_Float1718Output_2213);

SumNode_Float495: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1718Output_2213,ProductNode_Float1432Output_1845,SumNode_Float495Output_2214);

ProductNode_Float1719: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v6,SumNode_Float495Output_2214,ProductNode_Float1719Output_2215);

ProductNode_Float1720: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1720weight,v4,ProductNode_Float1720Output_2216);

ProductNode_Float1721: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1721weight,v8,ProductNode_Float1721Output_2217);

ProductNode_Float1722: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1722weight,vb8,ProductNode_Float1722Output_2218);

SumNode_Float496: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2Output_2,ProductNode_Float1Output_1,SumNode_Float496Output_2219);

ProductNode_Float1723: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v7,SumNode_Float0Output_3,ProductNode_Float1723Output_2220);

ProductNode_Float1724: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1724weight,v3,ProductNode_Float1724Output_2221);

ProductNode_Float1725: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1725weight,ProductNode_Float4Output_5,ProductNode_Float1725Output_2222);

ProductNode_Float1726: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1726weight,ProductNode_Float5Output_6,ProductNode_Float1726Output_2223);

ProductNode_Float1727: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1727weight,vb3,ProductNode_Float1727Output_2224);

ProductNode_Float1728: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1728weight,ProductNode_Float7Output_8,ProductNode_Float1728Output_2225);

ProductNode_Float1729: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1729weight,ProductNode_Float8Output_9,ProductNode_Float1729Output_2226);

SumNode_Float497: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float9Output_10,ProductNode_Float6Output_7,SumNode_Float497Output_2227);

ProductNode_Float1730: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float1Output_11,ProductNode_Float3Output_4,ProductNode_Float1730Output_2228);

ProductNode_Float1731: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1731weight,ProductNode_Float10Output_12,ProductNode_Float1731Output_2229);

ProductNode_Float1732: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1732weight,v8,ProductNode_Float1732Output_2230);

ProductNode_Float1733: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1733weight,vb8,ProductNode_Float1733Output_2231);

SumNode_Float498: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float13Output_15,ProductNode_Float12Output_14,SumNode_Float498Output_2232);

ProductNode_Float1734: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb7,SumNode_Float2Output_16,ProductNode_Float1734Output_2233);

ProductNode_Float1735: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1735weight,v3,ProductNode_Float1735Output_2234);

ProductNode_Float1736: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1736weight,ProductNode_Float4Output_5,ProductNode_Float1736Output_2235);

ProductNode_Float1737: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1737weight,ProductNode_Float16Output_19,ProductNode_Float1737Output_2236);

ProductNode_Float1738: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1738weight,vb3,ProductNode_Float1738Output_2237);

ProductNode_Float1739: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1739weight,ProductNode_Float7Output_8,ProductNode_Float1739Output_2238);

ProductNode_Float1740: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1740weight,ProductNode_Float19Output_22,ProductNode_Float1740Output_2239);

SumNode_Float499: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float20Output_23,ProductNode_Float17Output_20,SumNode_Float499Output_2240);

ProductNode_Float1741: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float3Output_24,ProductNode_Float14Output_17,ProductNode_Float1741Output_2241);

ProductNode_Float1742: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1742weight,ProductNode_Float21Output_25,ProductNode_Float1742Output_2242);

SumNode_Float500: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float595Output_764,ProductNode_Float584Output_751,SumNode_Float500Output_2243);

ProductNode_Float1743: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float169Output_765,ProductNode_Float0Output_0,ProductNode_Float1743Output_2244);

ProductNode_Float1744: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1744weight,ProductNode_Float596Output_766,ProductNode_Float1744Output_2245);

ProductNode_Float1745: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1745weight,vb4,ProductNode_Float1745Output_2246);

ProductNode_Float1746: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1746weight,v8,ProductNode_Float1746Output_2247);

ProductNode_Float1747: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1747weight,vb8,ProductNode_Float1747Output_2248);

SumNode_Float501: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float27Output_32,ProductNode_Float26Output_31,SumNode_Float501Output_2249);

ProductNode_Float1748: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v7,SumNode_Float5Output_33,ProductNode_Float1748Output_2250);

ProductNode_Float1749: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1749weight,v3,ProductNode_Float1749Output_2251);

ProductNode_Float1750: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1750weight,ProductNode_Float29Output_35,ProductNode_Float1750Output_2252);

ProductNode_Float1751: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1751weight,ProductNode_Float30Output_36,ProductNode_Float1751Output_2253);

ProductNode_Float1752: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1752weight,vb3,ProductNode_Float1752Output_2254);

ProductNode_Float1753: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1753weight,ProductNode_Float32Output_38,ProductNode_Float1753Output_2255);

ProductNode_Float1754: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1754weight,ProductNode_Float33Output_39,ProductNode_Float1754Output_2256);

SumNode_Float502: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float34Output_40,ProductNode_Float31Output_37,SumNode_Float502Output_2257);

ProductNode_Float1755: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float6Output_41,ProductNode_Float28Output_34,ProductNode_Float1755Output_2258);

ProductNode_Float1756: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1756weight,ProductNode_Float35Output_42,ProductNode_Float1756Output_2259);

ProductNode_Float1757: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1757weight,v8,ProductNode_Float1757Output_2260);

ProductNode_Float1758: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1758weight,vb8,ProductNode_Float1758Output_2261);

SumNode_Float503: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float38Output_45,ProductNode_Float37Output_44,SumNode_Float503Output_2262);

ProductNode_Float1759: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb7,SumNode_Float7Output_46,ProductNode_Float1759Output_2263);

ProductNode_Float1760: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1760weight,v3,ProductNode_Float1760Output_2264);

ProductNode_Float1761: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1761weight,ProductNode_Float29Output_35,ProductNode_Float1761Output_2265);

ProductNode_Float1762: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1762weight,ProductNode_Float41Output_49,ProductNode_Float1762Output_2266);

ProductNode_Float1763: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1763weight,vb3,ProductNode_Float1763Output_2267);

ProductNode_Float1764: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1764weight,ProductNode_Float32Output_38,ProductNode_Float1764Output_2268);

ProductNode_Float1765: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1765weight,ProductNode_Float44Output_52,ProductNode_Float1765Output_2269);

SumNode_Float504: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float45Output_53,ProductNode_Float42Output_50,SumNode_Float504Output_2270);

ProductNode_Float1766: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float8Output_54,ProductNode_Float39Output_47,ProductNode_Float1766Output_2271);

ProductNode_Float1767: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1767weight,ProductNode_Float46Output_55,ProductNode_Float1767Output_2272);

SumNode_Float505: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float620Output_794,ProductNode_Float609Output_781,SumNode_Float505Output_2273);

ProductNode_Float1768: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float174Output_795,ProductNode_Float25Output_30,ProductNode_Float1768Output_2274);

ProductNode_Float1769: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1769weight,ProductNode_Float621Output_796,ProductNode_Float1769Output_2275);

SumNode_Float506: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float622Output_797,ProductNode_Float597Output_767,SumNode_Float506Output_2276);

ProductNode_Float1770: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v5,SumNode_Float175Output_798,ProductNode_Float1770Output_2277);

ProductNode_Float1771: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1771weight,ProductNode_Float623Output_799,ProductNode_Float1771Output_2278);

ProductNode_Float1772: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1772weight,v4,ProductNode_Float1772Output_2279);

ProductNode_Float1773: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1773weight,v8,ProductNode_Float1773Output_2280);

ProductNode_Float1774: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1774weight,vb8,ProductNode_Float1774Output_2281);

SumNode_Float507: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float54Output_65,ProductNode_Float53Output_64,SumNode_Float507Output_2282);

ProductNode_Float1775: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v7,SumNode_Float11Output_66,ProductNode_Float1775Output_2283);

ProductNode_Float1776: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1776weight,v3,ProductNode_Float1776Output_2284);

ProductNode_Float1777: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1777weight,ProductNode_Float4Output_5,ProductNode_Float1777Output_2285);

ProductNode_Float1778: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1778weight,ProductNode_Float5Output_6,ProductNode_Float1778Output_2286);

ProductNode_Float1779: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1779weight,vb3,ProductNode_Float1779Output_2287);

ProductNode_Float1780: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1780weight,ProductNode_Float7Output_8,ProductNode_Float1780Output_2288);

ProductNode_Float1781: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1781weight,ProductNode_Float8Output_9,ProductNode_Float1781Output_2289);

SumNode_Float508: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float61Output_73,ProductNode_Float58Output_70,SumNode_Float508Output_2290);

ProductNode_Float1782: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float12Output_74,ProductNode_Float55Output_67,ProductNode_Float1782Output_2291);

ProductNode_Float1783: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1783weight,ProductNode_Float62Output_75,ProductNode_Float1783Output_2292);

ProductNode_Float1784: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1784weight,v8,ProductNode_Float1784Output_2293);

ProductNode_Float1785: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1785weight,vb8,ProductNode_Float1785Output_2294);

SumNode_Float509: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float65Output_78,ProductNode_Float64Output_77,SumNode_Float509Output_2295);

ProductNode_Float1786: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb7,SumNode_Float13Output_79,ProductNode_Float1786Output_2296);

ProductNode_Float1787: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1787weight,v3,ProductNode_Float1787Output_2297);

ProductNode_Float1788: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1788weight,ProductNode_Float4Output_5,ProductNode_Float1788Output_2298);

ProductNode_Float1789: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1789weight,ProductNode_Float16Output_19,ProductNode_Float1789Output_2299);

ProductNode_Float1790: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1790weight,vb3,ProductNode_Float1790Output_2300);

ProductNode_Float1791: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1791weight,ProductNode_Float7Output_8,ProductNode_Float1791Output_2301);

ProductNode_Float1792: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1792weight,ProductNode_Float19Output_22,ProductNode_Float1792Output_2302);

SumNode_Float510: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float72Output_86,ProductNode_Float69Output_83,SumNode_Float510Output_2303);

ProductNode_Float1793: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float14Output_87,ProductNode_Float66Output_80,ProductNode_Float1793Output_2304);

ProductNode_Float1794: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1794weight,ProductNode_Float73Output_88,ProductNode_Float1794Output_2305);

SumNode_Float511: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float647Output_827,ProductNode_Float636Output_814,SumNode_Float511Output_2306);

ProductNode_Float1795: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float180Output_828,ProductNode_Float0Output_0,ProductNode_Float1795Output_2307);

ProductNode_Float1796: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1796weight,ProductNode_Float648Output_829,ProductNode_Float1796Output_2308);

ProductNode_Float1797: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1797weight,vb4,ProductNode_Float1797Output_2309);

ProductNode_Float1798: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1798weight,v8,ProductNode_Float1798Output_2310);

ProductNode_Float1799: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1799weight,vb8,ProductNode_Float1799Output_2311);

SumNode_Float512: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float79Output_95,ProductNode_Float78Output_94,SumNode_Float512Output_2312);

ProductNode_Float1800: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v7,SumNode_Float16Output_96,ProductNode_Float1800Output_2313);

ProductNode_Float1801: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1801weight,v3,ProductNode_Float1801Output_2314);

ProductNode_Float1802: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1802weight,ProductNode_Float29Output_35,ProductNode_Float1802Output_2315);

ProductNode_Float1803: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1803weight,ProductNode_Float30Output_36,ProductNode_Float1803Output_2316);

ProductNode_Float1804: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1804weight,vb3,ProductNode_Float1804Output_2317);

ProductNode_Float1805: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1805weight,ProductNode_Float32Output_38,ProductNode_Float1805Output_2318);

ProductNode_Float1806: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1806weight,ProductNode_Float33Output_39,ProductNode_Float1806Output_2319);

SumNode_Float513: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float86Output_103,ProductNode_Float83Output_100,SumNode_Float513Output_2320);

ProductNode_Float1807: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float17Output_104,ProductNode_Float80Output_97,ProductNode_Float1807Output_2321);

ProductNode_Float1808: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1808weight,ProductNode_Float87Output_105,ProductNode_Float1808Output_2322);

ProductNode_Float1809: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1809weight,v8,ProductNode_Float1809Output_2323);

ProductNode_Float1810: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1810weight,vb8,ProductNode_Float1810Output_2324);

SumNode_Float514: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float90Output_108,ProductNode_Float89Output_107,SumNode_Float514Output_2325);

ProductNode_Float1811: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb7,SumNode_Float18Output_109,ProductNode_Float1811Output_2326);

ProductNode_Float1812: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1812weight,v3,ProductNode_Float1812Output_2327);

ProductNode_Float1813: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1813weight,ProductNode_Float29Output_35,ProductNode_Float1813Output_2328);

ProductNode_Float1814: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1814weight,ProductNode_Float41Output_49,ProductNode_Float1814Output_2329);

ProductNode_Float1815: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1815weight,vb3,ProductNode_Float1815Output_2330);

ProductNode_Float1816: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1816weight,ProductNode_Float32Output_38,ProductNode_Float1816Output_2331);

ProductNode_Float1817: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1817weight,ProductNode_Float44Output_52,ProductNode_Float1817Output_2332);

SumNode_Float515: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float97Output_116,ProductNode_Float94Output_113,SumNode_Float515Output_2333);

ProductNode_Float1818: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float19Output_117,ProductNode_Float91Output_110,ProductNode_Float1818Output_2334);

ProductNode_Float1819: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1819weight,ProductNode_Float98Output_118,ProductNode_Float1819Output_2335);

SumNode_Float516: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float672Output_857,ProductNode_Float661Output_844,SumNode_Float516Output_2336);

ProductNode_Float1820: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float185Output_858,ProductNode_Float25Output_30,ProductNode_Float1820Output_2337);

ProductNode_Float1821: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1821weight,ProductNode_Float673Output_859,ProductNode_Float1821Output_2338);

SumNode_Float517: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float674Output_860,ProductNode_Float649Output_830,SumNode_Float517Output_2339);

ProductNode_Float1822: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb5,SumNode_Float186Output_861,ProductNode_Float1822Output_2340);

ProductNode_Float1823: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1823weight,ProductNode_Float675Output_862,ProductNode_Float1823Output_2341);

SumNode_Float518: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1823Output_2341,ProductNode_Float1771Output_2278,SumNode_Float518Output_2342);

ProductNode_Float1824: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v16,SumNode_Float518Output_2342,ProductNode_Float1824Output_2343);

ProductNode_Float1825: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1825weight,v11,ProductNode_Float1825Output_2344);

ProductNode_Float1826: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1826weight,vb11,ProductNode_Float1826Output_2345);

SumNode_Float519: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float679Output_867,ProductNode_Float678Output_866,SumNode_Float519Output_2346);

ProductNode_Float1827: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v12,SumNode_Float188Output_868,ProductNode_Float1827Output_2347);

ProductNode_Float1828: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1828weight,ProductNode_Float680Output_869,ProductNode_Float1828Output_2348);

ProductNode_Float1829: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1829weight,v2,ProductNode_Float1829Output_2349);

ProductNode_Float1830: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1830weight,vb2,ProductNode_Float1830Output_2350);

SumNode_Float520: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float110Output_134,ProductNode_Float109Output_133,SumNode_Float520Output_2351);

ProductNode_Float1831: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float24Output_135,ProductNode_Float681Output_870,ProductNode_Float1831Output_2352);

ProductNode_Float1832: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1832weight,v11,ProductNode_Float1832Output_2353);

ProductNode_Float1833: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1833weight,vb11,ProductNode_Float1833Output_2354);

SumNode_Float521: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float686Output_876,ProductNode_Float685Output_875,SumNode_Float521Output_2355);

ProductNode_Float1834: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb12,SumNode_Float190Output_877,ProductNode_Float1834Output_2356);

ProductNode_Float1835: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1835weight,ProductNode_Float687Output_878,ProductNode_Float1835Output_2357);

ProductNode_Float1836: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1836weight,v2,ProductNode_Float1836Output_2358);

ProductNode_Float1837: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1837weight,vb2,ProductNode_Float1837Output_2359);

SumNode_Float522: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float117Output_143,ProductNode_Float116Output_142,SumNode_Float522Output_2360);

ProductNode_Float1838: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float26Output_144,ProductNode_Float688Output_879,ProductNode_Float1838Output_2361);

SumNode_Float523: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float691Output_883,ProductNode_Float684Output_874,SumNode_Float523Output_2362);

ProductNode_Float1839: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v13,SumNode_Float192Output_884,ProductNode_Float1839Output_2363);

ProductNode_Float1840: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1840weight,ProductNode_Float692Output_885,ProductNode_Float1840Output_2364);

ProductNode_Float1841: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1841weight,v11,ProductNode_Float1841Output_2365);

ProductNode_Float1842: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1842weight,vb11,ProductNode_Float1842Output_2366);

SumNode_Float524: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float695Output_888,ProductNode_Float694Output_887,SumNode_Float524Output_2367);

ProductNode_Float1843: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v12,SumNode_Float193Output_889,ProductNode_Float1843Output_2368);

ProductNode_Float1844: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1844weight,ProductNode_Float696Output_890,ProductNode_Float1844Output_2369);

ProductNode_Float1845: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1845weight,v2,ProductNode_Float1845Output_2370);

ProductNode_Float1846: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1846weight,vb2,ProductNode_Float1846Output_2371);

SumNode_Float525: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float126Output_155,ProductNode_Float125Output_154,SumNode_Float525Output_2372);

ProductNode_Float1847: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float29Output_156,ProductNode_Float697Output_891,ProductNode_Float1847Output_2373);

ProductNode_Float1848: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1848weight,v11,ProductNode_Float1848Output_2374);

ProductNode_Float1849: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1849weight,vb11,ProductNode_Float1849Output_2375);

SumNode_Float526: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float702Output_897,ProductNode_Float701Output_896,SumNode_Float526Output_2376);

ProductNode_Float1850: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb12,SumNode_Float195Output_898,ProductNode_Float1850Output_2377);

ProductNode_Float1851: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1851weight,ProductNode_Float703Output_899,ProductNode_Float1851Output_2378);

ProductNode_Float1852: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1852weight,v2,ProductNode_Float1852Output_2379);

ProductNode_Float1853: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1853weight,vb2,ProductNode_Float1853Output_2380);

SumNode_Float527: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float133Output_164,ProductNode_Float132Output_163,SumNode_Float527Output_2381);

ProductNode_Float1854: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float31Output_165,ProductNode_Float704Output_900,ProductNode_Float1854Output_2382);

SumNode_Float528: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float707Output_904,ProductNode_Float700Output_895,SumNode_Float528Output_2383);

ProductNode_Float1855: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb13,SumNode_Float197Output_905,ProductNode_Float1855Output_2384);

ProductNode_Float1856: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1856weight,ProductNode_Float708Output_906,ProductNode_Float1856Output_2385);

SumNode_Float529: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float709Output_907,ProductNode_Float693Output_886,SumNode_Float529Output_2386);

ProductNode_Float1857: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v10,SumNode_Float198Output_908,ProductNode_Float1857Output_2387);

ProductNode_Float1858: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1858weight,v1,ProductNode_Float1858Output_2388);

ProductNode_Float1859: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1859weight,vb1,ProductNode_Float1859Output_2389);

SumNode_Float530: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1286Output_1651,ProductNode_Float1285Output_1650,SumNode_Float530Output_2390);

ProductNode_Float1860: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v9,SumNode_Float365Output_1652,ProductNode_Float1860Output_2391);

ProductNode_Float1861: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1861weight,ProductNode_Float1287Output_1653,ProductNode_Float1861Output_2392);

ProductNode_Float1862: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1862weight,ProductNode_Float1288Output_1654,ProductNode_Float1862Output_2393);

ProductNode_Float1863: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1863weight,v1,ProductNode_Float1863Output_2394);

ProductNode_Float1864: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1864weight,vb1,ProductNode_Float1864Output_2395);

SumNode_Float531: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1291Output_1657,ProductNode_Float1290Output_1656,SumNode_Float531Output_2396);

ProductNode_Float1865: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb9,SumNode_Float366Output_1658,ProductNode_Float1865Output_2397);

ProductNode_Float1866: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1866weight,ProductNode_Float1292Output_1659,ProductNode_Float1866Output_2398);

ProductNode_Float1867: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1867weight,ProductNode_Float1293Output_1660,ProductNode_Float1867Output_2399);

SumNode_Float532: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1294Output_1661,ProductNode_Float1289Output_1655,SumNode_Float532Output_2400);

ProductNode_Float1868: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float367Output_1662,ProductNode_Float710Output_909,ProductNode_Float1868Output_2401);

ProductNode_Float1869: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1869weight,v11,ProductNode_Float1869Output_2402);

ProductNode_Float1870: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1870weight,vb11,ProductNode_Float1870Output_2403);

SumNode_Float533: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float679Output_867,ProductNode_Float678Output_866,SumNode_Float533Output_2404);

ProductNode_Float1871: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v12,SumNode_Float188Output_868,ProductNode_Float1871Output_2405);

ProductNode_Float1872: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1872weight,ProductNode_Float680Output_869,ProductNode_Float1872Output_2406);

ProductNode_Float1873: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1873weight,v2,ProductNode_Float1873Output_2407);

ProductNode_Float1874: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1874weight,vb2,ProductNode_Float1874Output_2408);

SumNode_Float534: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float110Output_134,ProductNode_Float109Output_133,SumNode_Float534Output_2409);

ProductNode_Float1875: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float24Output_135,ProductNode_Float681Output_870,ProductNode_Float1875Output_2410);

ProductNode_Float1876: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1876weight,v11,ProductNode_Float1876Output_2411);

ProductNode_Float1877: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1877weight,vb11,ProductNode_Float1877Output_2412);

SumNode_Float535: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float686Output_876,ProductNode_Float685Output_875,SumNode_Float535Output_2413);

ProductNode_Float1878: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb12,SumNode_Float190Output_877,ProductNode_Float1878Output_2414);

ProductNode_Float1879: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1879weight,ProductNode_Float687Output_878,ProductNode_Float1879Output_2415);

ProductNode_Float1880: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1880weight,v2,ProductNode_Float1880Output_2416);

ProductNode_Float1881: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1881weight,vb2,ProductNode_Float1881Output_2417);

SumNode_Float536: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float117Output_143,ProductNode_Float116Output_142,SumNode_Float536Output_2418);

ProductNode_Float1882: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float26Output_144,ProductNode_Float688Output_879,ProductNode_Float1882Output_2419);

SumNode_Float537: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float691Output_883,ProductNode_Float684Output_874,SumNode_Float537Output_2420);

ProductNode_Float1883: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v13,SumNode_Float192Output_884,ProductNode_Float1883Output_2421);

ProductNode_Float1884: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1884weight,ProductNode_Float692Output_885,ProductNode_Float1884Output_2422);

ProductNode_Float1885: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1885weight,v11,ProductNode_Float1885Output_2423);

ProductNode_Float1886: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1886weight,vb11,ProductNode_Float1886Output_2424);

SumNode_Float538: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float695Output_888,ProductNode_Float694Output_887,SumNode_Float538Output_2425);

ProductNode_Float1887: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v12,SumNode_Float193Output_889,ProductNode_Float1887Output_2426);

ProductNode_Float1888: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1888weight,ProductNode_Float696Output_890,ProductNode_Float1888Output_2427);

ProductNode_Float1889: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1889weight,v2,ProductNode_Float1889Output_2428);

ProductNode_Float1890: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1890weight,vb2,ProductNode_Float1890Output_2429);

SumNode_Float539: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float126Output_155,ProductNode_Float125Output_154,SumNode_Float539Output_2430);

ProductNode_Float1891: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float29Output_156,ProductNode_Float697Output_891,ProductNode_Float1891Output_2431);

ProductNode_Float1892: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1892weight,v11,ProductNode_Float1892Output_2432);

ProductNode_Float1893: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1893weight,vb11,ProductNode_Float1893Output_2433);

SumNode_Float540: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float702Output_897,ProductNode_Float701Output_896,SumNode_Float540Output_2434);

ProductNode_Float1894: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb12,SumNode_Float195Output_898,ProductNode_Float1894Output_2435);

ProductNode_Float1895: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1895weight,ProductNode_Float703Output_899,ProductNode_Float1895Output_2436);

ProductNode_Float1896: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1896weight,v2,ProductNode_Float1896Output_2437);

ProductNode_Float1897: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1897weight,vb2,ProductNode_Float1897Output_2438);

SumNode_Float541: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float133Output_164,ProductNode_Float132Output_163,SumNode_Float541Output_2439);

ProductNode_Float1898: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float31Output_165,ProductNode_Float704Output_900,ProductNode_Float1898Output_2440);

SumNode_Float542: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float707Output_904,ProductNode_Float700Output_895,SumNode_Float542Output_2441);

ProductNode_Float1899: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb13,SumNode_Float197Output_905,ProductNode_Float1899Output_2442);

ProductNode_Float1900: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1900weight,ProductNode_Float708Output_906,ProductNode_Float1900Output_2443);

SumNode_Float543: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float753Output_965,ProductNode_Float737Output_944,SumNode_Float543Output_2444);

ProductNode_Float1901: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb10,SumNode_Float212Output_966,ProductNode_Float1901Output_2445);

ProductNode_Float1902: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1902weight,v1,ProductNode_Float1902Output_2446);

ProductNode_Float1903: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1903weight,vb1,ProductNode_Float1903Output_2447);

SumNode_Float544: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1330Output_1709,ProductNode_Float1329Output_1708,SumNode_Float544Output_2448);

ProductNode_Float1904: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v9,SumNode_Float379Output_1710,ProductNode_Float1904Output_2449);

ProductNode_Float1905: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1905weight,ProductNode_Float1331Output_1711,ProductNode_Float1905Output_2450);

ProductNode_Float1906: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1906weight,ProductNode_Float1332Output_1712,ProductNode_Float1906Output_2451);

ProductNode_Float1907: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1907weight,v1,ProductNode_Float1907Output_2452);

ProductNode_Float1908: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1908weight,vb1,ProductNode_Float1908Output_2453);

SumNode_Float545: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1335Output_1715,ProductNode_Float1334Output_1714,SumNode_Float545Output_2454);

ProductNode_Float1909: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb9,SumNode_Float380Output_1716,ProductNode_Float1909Output_2455);

ProductNode_Float1910: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1910weight,ProductNode_Float1336Output_1717,ProductNode_Float1910Output_2456);

ProductNode_Float1911: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1911weight,ProductNode_Float1337Output_1718,ProductNode_Float1911Output_2457);

SumNode_Float546: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1338Output_1719,ProductNode_Float1333Output_1713,SumNode_Float546Output_2458);

ProductNode_Float1912: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float381Output_1720,ProductNode_Float754Output_967,ProductNode_Float1912Output_2459);

SumNode_Float547: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1912Output_2459,ProductNode_Float1868Output_2401,SumNode_Float547Output_2460);

ProductNode_Float1913: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v15,SumNode_Float547Output_2460,ProductNode_Float1913Output_2461);

ProductNode_Float1914: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1914weight,ProductNode_Float1913Output_2461,ProductNode_Float1914Output_2462);

ProductNode_Float1915: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1915weight,v11,ProductNode_Float1915Output_2463);

ProductNode_Float1916: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1916weight,vb11,ProductNode_Float1916Output_2464);

SumNode_Float548: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float679Output_867,ProductNode_Float678Output_866,SumNode_Float548Output_2465);

ProductNode_Float1917: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v12,SumNode_Float188Output_868,ProductNode_Float1917Output_2466);

ProductNode_Float1918: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1918weight,ProductNode_Float680Output_869,ProductNode_Float1918Output_2467);

ProductNode_Float1919: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1919weight,v2,ProductNode_Float1919Output_2468);

ProductNode_Float1920: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1920weight,vb2,ProductNode_Float1920Output_2469);

SumNode_Float549: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float200Output_253,ProductNode_Float199Output_252,SumNode_Float549Output_2470);

ProductNode_Float1921: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float53Output_254,ProductNode_Float681Output_870,ProductNode_Float1921Output_2471);

ProductNode_Float1922: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1922weight,v11,ProductNode_Float1922Output_2472);

ProductNode_Float1923: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1923weight,vb11,ProductNode_Float1923Output_2473);

SumNode_Float550: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float686Output_876,ProductNode_Float685Output_875,SumNode_Float550Output_2474);

ProductNode_Float1924: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb12,SumNode_Float190Output_877,ProductNode_Float1924Output_2475);

ProductNode_Float1925: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1925weight,ProductNode_Float687Output_878,ProductNode_Float1925Output_2476);

ProductNode_Float1926: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1926weight,v2,ProductNode_Float1926Output_2477);

ProductNode_Float1927: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1927weight,vb2,ProductNode_Float1927Output_2478);

SumNode_Float551: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float207Output_262,ProductNode_Float206Output_261,SumNode_Float551Output_2479);

ProductNode_Float1928: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float55Output_263,ProductNode_Float688Output_879,ProductNode_Float1928Output_2480);

SumNode_Float552: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float781Output_1002,ProductNode_Float774Output_993,SumNode_Float552Output_2481);

ProductNode_Float1929: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v13,SumNode_Float221Output_1003,ProductNode_Float1929Output_2482);

ProductNode_Float1930: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1930weight,ProductNode_Float782Output_1004,ProductNode_Float1930Output_2483);

ProductNode_Float1931: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1931weight,v11,ProductNode_Float1931Output_2484);

ProductNode_Float1932: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1932weight,vb11,ProductNode_Float1932Output_2485);

SumNode_Float553: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float695Output_888,ProductNode_Float694Output_887,SumNode_Float553Output_2486);

ProductNode_Float1933: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v12,SumNode_Float193Output_889,ProductNode_Float1933Output_2487);

ProductNode_Float1934: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1934weight,ProductNode_Float696Output_890,ProductNode_Float1934Output_2488);

ProductNode_Float1935: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1935weight,v2,ProductNode_Float1935Output_2489);

ProductNode_Float1936: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1936weight,vb2,ProductNode_Float1936Output_2490);

SumNode_Float554: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float216Output_274,ProductNode_Float215Output_273,SumNode_Float554Output_2491);

ProductNode_Float1937: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float58Output_275,ProductNode_Float697Output_891,ProductNode_Float1937Output_2492);

ProductNode_Float1938: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1938weight,v11,ProductNode_Float1938Output_2493);

ProductNode_Float1939: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1939weight,vb11,ProductNode_Float1939Output_2494);

SumNode_Float555: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float702Output_897,ProductNode_Float701Output_896,SumNode_Float555Output_2495);

ProductNode_Float1940: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb12,SumNode_Float195Output_898,ProductNode_Float1940Output_2496);

ProductNode_Float1941: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1941weight,ProductNode_Float703Output_899,ProductNode_Float1941Output_2497);

ProductNode_Float1942: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1942weight,v2,ProductNode_Float1942Output_2498);

ProductNode_Float1943: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1943weight,vb2,ProductNode_Float1943Output_2499);

SumNode_Float556: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float223Output_283,ProductNode_Float222Output_282,SumNode_Float556Output_2500);

ProductNode_Float1944: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float60Output_284,ProductNode_Float704Output_900,ProductNode_Float1944Output_2501);

SumNode_Float557: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float797Output_1023,ProductNode_Float790Output_1014,SumNode_Float557Output_2502);

ProductNode_Float1945: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb13,SumNode_Float226Output_1024,ProductNode_Float1945Output_2503);

ProductNode_Float1946: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1946weight,ProductNode_Float798Output_1025,ProductNode_Float1946Output_2504);

SumNode_Float558: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float799Output_1026,ProductNode_Float783Output_1005,SumNode_Float558Output_2505);

ProductNode_Float1947: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v10,SumNode_Float227Output_1027,ProductNode_Float1947Output_2506);

ProductNode_Float1948: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1948weight,v1,ProductNode_Float1948Output_2507);

ProductNode_Float1949: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1949weight,vb1,ProductNode_Float1949Output_2508);

SumNode_Float559: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1286Output_1651,ProductNode_Float1285Output_1650,SumNode_Float559Output_2509);

ProductNode_Float1950: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v9,SumNode_Float365Output_1652,ProductNode_Float1950Output_2510);

ProductNode_Float1951: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1951weight,ProductNode_Float1287Output_1653,ProductNode_Float1951Output_2511);

ProductNode_Float1952: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1952weight,ProductNode_Float1378Output_1773,ProductNode_Float1952Output_2512);

ProductNode_Float1953: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1953weight,v1,ProductNode_Float1953Output_2513);

ProductNode_Float1954: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1954weight,vb1,ProductNode_Float1954Output_2514);

SumNode_Float560: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1291Output_1657,ProductNode_Float1290Output_1656,SumNode_Float560Output_2515);

ProductNode_Float1955: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb9,SumNode_Float366Output_1658,ProductNode_Float1955Output_2516);

ProductNode_Float1956: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1956weight,ProductNode_Float1292Output_1659,ProductNode_Float1956Output_2517);

ProductNode_Float1957: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1957weight,ProductNode_Float1383Output_1779,ProductNode_Float1957Output_2518);

SumNode_Float561: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1384Output_1780,ProductNode_Float1379Output_1774,SumNode_Float561Output_2519);

ProductNode_Float1958: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float396Output_1781,ProductNode_Float800Output_1028,ProductNode_Float1958Output_2520);

ProductNode_Float1959: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1959weight,v11,ProductNode_Float1959Output_2521);

ProductNode_Float1960: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1960weight,vb11,ProductNode_Float1960Output_2522);

SumNode_Float562: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float679Output_867,ProductNode_Float678Output_866,SumNode_Float562Output_2523);

ProductNode_Float1961: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v12,SumNode_Float188Output_868,ProductNode_Float1961Output_2524);

ProductNode_Float1962: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1962weight,ProductNode_Float680Output_869,ProductNode_Float1962Output_2525);

ProductNode_Float1963: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1963weight,v2,ProductNode_Float1963Output_2526);

ProductNode_Float1964: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1964weight,vb2,ProductNode_Float1964Output_2527);

SumNode_Float563: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float200Output_253,ProductNode_Float199Output_252,SumNode_Float563Output_2528);

ProductNode_Float1965: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float53Output_254,ProductNode_Float681Output_870,ProductNode_Float1965Output_2529);

ProductNode_Float1966: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1966weight,v11,ProductNode_Float1966Output_2530);

ProductNode_Float1967: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1967weight,vb11,ProductNode_Float1967Output_2531);

SumNode_Float564: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float686Output_876,ProductNode_Float685Output_875,SumNode_Float564Output_2532);

ProductNode_Float1968: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb12,SumNode_Float190Output_877,ProductNode_Float1968Output_2533);

ProductNode_Float1969: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1969weight,ProductNode_Float687Output_878,ProductNode_Float1969Output_2534);

ProductNode_Float1970: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1970weight,v2,ProductNode_Float1970Output_2535);

ProductNode_Float1971: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1971weight,vb2,ProductNode_Float1971Output_2536);

SumNode_Float565: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float207Output_262,ProductNode_Float206Output_261,SumNode_Float565Output_2537);

ProductNode_Float1972: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float55Output_263,ProductNode_Float688Output_879,ProductNode_Float1972Output_2538);

SumNode_Float566: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float781Output_1002,ProductNode_Float774Output_993,SumNode_Float566Output_2539);

ProductNode_Float1973: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v13,SumNode_Float221Output_1003,ProductNode_Float1973Output_2540);

ProductNode_Float1974: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1974weight,ProductNode_Float782Output_1004,ProductNode_Float1974Output_2541);

ProductNode_Float1975: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1975weight,v11,ProductNode_Float1975Output_2542);

ProductNode_Float1976: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1976weight,vb11,ProductNode_Float1976Output_2543);

SumNode_Float567: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float695Output_888,ProductNode_Float694Output_887,SumNode_Float567Output_2544);

ProductNode_Float1977: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v12,SumNode_Float193Output_889,ProductNode_Float1977Output_2545);

ProductNode_Float1978: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1978weight,ProductNode_Float696Output_890,ProductNode_Float1978Output_2546);

ProductNode_Float1979: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1979weight,v2,ProductNode_Float1979Output_2547);

ProductNode_Float1980: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1980weight,vb2,ProductNode_Float1980Output_2548);

SumNode_Float568: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float216Output_274,ProductNode_Float215Output_273,SumNode_Float568Output_2549);

ProductNode_Float1981: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float58Output_275,ProductNode_Float697Output_891,ProductNode_Float1981Output_2550);

ProductNode_Float1982: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1982weight,v11,ProductNode_Float1982Output_2551);

ProductNode_Float1983: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1983weight,vb11,ProductNode_Float1983Output_2552);

SumNode_Float569: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float702Output_897,ProductNode_Float701Output_896,SumNode_Float569Output_2553);

ProductNode_Float1984: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb12,SumNode_Float195Output_898,ProductNode_Float1984Output_2554);

ProductNode_Float1985: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1985weight,ProductNode_Float703Output_899,ProductNode_Float1985Output_2555);

ProductNode_Float1986: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1986weight,v2,ProductNode_Float1986Output_2556);

ProductNode_Float1987: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1987weight,vb2,ProductNode_Float1987Output_2557);

SumNode_Float570: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float223Output_283,ProductNode_Float222Output_282,SumNode_Float570Output_2558);

ProductNode_Float1988: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float60Output_284,ProductNode_Float704Output_900,ProductNode_Float1988Output_2559);

SumNode_Float571: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float797Output_1023,ProductNode_Float790Output_1014,SumNode_Float571Output_2560);

ProductNode_Float1989: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb13,SumNode_Float226Output_1024,ProductNode_Float1989Output_2561);

ProductNode_Float1990: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1990weight,ProductNode_Float798Output_1025,ProductNode_Float1990Output_2562);

SumNode_Float572: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float843Output_1084,ProductNode_Float827Output_1063,SumNode_Float572Output_2563);

ProductNode_Float1991: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb10,SumNode_Float241Output_1085,ProductNode_Float1991Output_2564);

ProductNode_Float1992: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1992weight,v1,ProductNode_Float1992Output_2565);

ProductNode_Float1993: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1993weight,vb1,ProductNode_Float1993Output_2566);

SumNode_Float573: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1330Output_1709,ProductNode_Float1329Output_1708,SumNode_Float573Output_2567);

ProductNode_Float1994: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v9,SumNode_Float379Output_1710,ProductNode_Float1994Output_2568);

ProductNode_Float1995: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1995weight,ProductNode_Float1331Output_1711,ProductNode_Float1995Output_2569);

ProductNode_Float1996: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1996weight,ProductNode_Float1422Output_1831,ProductNode_Float1996Output_2570);

ProductNode_Float1997: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1997weight,v1,ProductNode_Float1997Output_2571);

ProductNode_Float1998: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1998weight,vb1,ProductNode_Float1998Output_2572);

SumNode_Float574: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1335Output_1715,ProductNode_Float1334Output_1714,SumNode_Float574Output_2573);

ProductNode_Float1999: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb9,SumNode_Float380Output_1716,ProductNode_Float1999Output_2574);

ProductNode_Float2000: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2000weight,ProductNode_Float1336Output_1717,ProductNode_Float2000Output_2575);

ProductNode_Float2001: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2001weight,ProductNode_Float1427Output_1837,ProductNode_Float2001Output_2576);

SumNode_Float575: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1428Output_1838,ProductNode_Float1423Output_1832,SumNode_Float575Output_2577);

ProductNode_Float2002: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float410Output_1839,ProductNode_Float844Output_1086,ProductNode_Float2002Output_2578);

SumNode_Float576: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2002Output_2578,ProductNode_Float1958Output_2520,SumNode_Float576Output_2579);

ProductNode_Float2003: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb15,SumNode_Float576Output_2579,ProductNode_Float2003Output_2580);

ProductNode_Float2004: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2004weight,ProductNode_Float2003Output_2580,ProductNode_Float2004Output_2581);

SumNode_Float577: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2004Output_2581,ProductNode_Float1914Output_2462,SumNode_Float577Output_2582);

ProductNode_Float2005: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float577Output_2582,ProductNode_Float1824Output_2343,ProductNode_Float2005Output_2583);

ProductNode_Float2006: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2006weight,v4,ProductNode_Float2006Output_2584);

ProductNode_Float2007: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2007weight,v8,ProductNode_Float2007Output_2585);

ProductNode_Float2008: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2008weight,vb8,ProductNode_Float2008Output_2586);

SumNode_Float578: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2Output_2,ProductNode_Float1Output_1,SumNode_Float578Output_2587);

ProductNode_Float2009: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v7,SumNode_Float0Output_3,ProductNode_Float2009Output_2588);

ProductNode_Float2010: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2010weight,v3,ProductNode_Float2010Output_2589);

ProductNode_Float2011: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2011weight,ProductNode_Float4Output_5,ProductNode_Float2011Output_2590);

ProductNode_Float2012: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2012weight,ProductNode_Float5Output_6,ProductNode_Float2012Output_2591);

ProductNode_Float2013: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2013weight,vb3,ProductNode_Float2013Output_2592);

ProductNode_Float2014: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2014weight,ProductNode_Float7Output_8,ProductNode_Float2014Output_2593);

ProductNode_Float2015: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2015weight,ProductNode_Float8Output_9,ProductNode_Float2015Output_2594);

SumNode_Float579: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float9Output_10,ProductNode_Float6Output_7,SumNode_Float579Output_2595);

ProductNode_Float2016: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float1Output_11,ProductNode_Float3Output_4,ProductNode_Float2016Output_2596);

ProductNode_Float2017: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2017weight,ProductNode_Float10Output_12,ProductNode_Float2017Output_2597);

ProductNode_Float2018: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2018weight,v8,ProductNode_Float2018Output_2598);

ProductNode_Float2019: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2019weight,vb8,ProductNode_Float2019Output_2599);

SumNode_Float580: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float13Output_15,ProductNode_Float12Output_14,SumNode_Float580Output_2600);

ProductNode_Float2020: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb7,SumNode_Float2Output_16,ProductNode_Float2020Output_2601);

ProductNode_Float2021: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2021weight,v3,ProductNode_Float2021Output_2602);

ProductNode_Float2022: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2022weight,ProductNode_Float4Output_5,ProductNode_Float2022Output_2603);

ProductNode_Float2023: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2023weight,ProductNode_Float16Output_19,ProductNode_Float2023Output_2604);

ProductNode_Float2024: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2024weight,vb3,ProductNode_Float2024Output_2605);

ProductNode_Float2025: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2025weight,ProductNode_Float7Output_8,ProductNode_Float2025Output_2606);

ProductNode_Float2026: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2026weight,ProductNode_Float19Output_22,ProductNode_Float2026Output_2607);

SumNode_Float581: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float20Output_23,ProductNode_Float17Output_20,SumNode_Float581Output_2608);

ProductNode_Float2027: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float3Output_24,ProductNode_Float14Output_17,ProductNode_Float2027Output_2609);

ProductNode_Float2028: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2028weight,ProductNode_Float21Output_25,ProductNode_Float2028Output_2610);

SumNode_Float582: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float595Output_764,ProductNode_Float584Output_751,SumNode_Float582Output_2611);

ProductNode_Float2029: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float169Output_765,ProductNode_Float0Output_0,ProductNode_Float2029Output_2612);

ProductNode_Float2030: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2030weight,ProductNode_Float596Output_766,ProductNode_Float2030Output_2613);

ProductNode_Float2031: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2031weight,vb4,ProductNode_Float2031Output_2614);

ProductNode_Float2032: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2032weight,v8,ProductNode_Float2032Output_2615);

ProductNode_Float2033: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2033weight,vb8,ProductNode_Float2033Output_2616);

SumNode_Float583: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float27Output_32,ProductNode_Float26Output_31,SumNode_Float583Output_2617);

ProductNode_Float2034: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v7,SumNode_Float5Output_33,ProductNode_Float2034Output_2618);

ProductNode_Float2035: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2035weight,v3,ProductNode_Float2035Output_2619);

ProductNode_Float2036: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2036weight,ProductNode_Float29Output_35,ProductNode_Float2036Output_2620);

ProductNode_Float2037: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2037weight,ProductNode_Float30Output_36,ProductNode_Float2037Output_2621);

ProductNode_Float2038: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2038weight,vb3,ProductNode_Float2038Output_2622);

ProductNode_Float2039: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2039weight,ProductNode_Float32Output_38,ProductNode_Float2039Output_2623);

ProductNode_Float2040: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2040weight,ProductNode_Float33Output_39,ProductNode_Float2040Output_2624);

SumNode_Float584: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float34Output_40,ProductNode_Float31Output_37,SumNode_Float584Output_2625);

ProductNode_Float2041: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float6Output_41,ProductNode_Float28Output_34,ProductNode_Float2041Output_2626);

ProductNode_Float2042: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2042weight,ProductNode_Float35Output_42,ProductNode_Float2042Output_2627);

ProductNode_Float2043: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2043weight,v8,ProductNode_Float2043Output_2628);

ProductNode_Float2044: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2044weight,vb8,ProductNode_Float2044Output_2629);

SumNode_Float585: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float38Output_45,ProductNode_Float37Output_44,SumNode_Float585Output_2630);

ProductNode_Float2045: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb7,SumNode_Float7Output_46,ProductNode_Float2045Output_2631);

ProductNode_Float2046: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2046weight,v3,ProductNode_Float2046Output_2632);

ProductNode_Float2047: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2047weight,ProductNode_Float29Output_35,ProductNode_Float2047Output_2633);

ProductNode_Float2048: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2048weight,ProductNode_Float41Output_49,ProductNode_Float2048Output_2634);

ProductNode_Float2049: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2049weight,vb3,ProductNode_Float2049Output_2635);

ProductNode_Float2050: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2050weight,ProductNode_Float32Output_38,ProductNode_Float2050Output_2636);

ProductNode_Float2051: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2051weight,ProductNode_Float44Output_52,ProductNode_Float2051Output_2637);

SumNode_Float586: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float45Output_53,ProductNode_Float42Output_50,SumNode_Float586Output_2638);

ProductNode_Float2052: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float8Output_54,ProductNode_Float39Output_47,ProductNode_Float2052Output_2639);

ProductNode_Float2053: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2053weight,ProductNode_Float46Output_55,ProductNode_Float2053Output_2640);

SumNode_Float587: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float620Output_794,ProductNode_Float609Output_781,SumNode_Float587Output_2641);

ProductNode_Float2054: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float174Output_795,ProductNode_Float25Output_30,ProductNode_Float2054Output_2642);

ProductNode_Float2055: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2055weight,ProductNode_Float621Output_796,ProductNode_Float2055Output_2643);

SumNode_Float588: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float908Output_1165,ProductNode_Float883Output_1135,SumNode_Float588Output_2644);

ProductNode_Float2056: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v5,SumNode_Float257Output_1166,ProductNode_Float2056Output_2645);

ProductNode_Float2057: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2057weight,ProductNode_Float909Output_1167,ProductNode_Float2057Output_2646);

ProductNode_Float2058: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2058weight,v4,ProductNode_Float2058Output_2647);

ProductNode_Float2059: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2059weight,v8,ProductNode_Float2059Output_2648);

ProductNode_Float2060: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2060weight,vb8,ProductNode_Float2060Output_2649);

SumNode_Float589: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float54Output_65,ProductNode_Float53Output_64,SumNode_Float589Output_2650);

ProductNode_Float2061: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v7,SumNode_Float11Output_66,ProductNode_Float2061Output_2651);

ProductNode_Float2062: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2062weight,v3,ProductNode_Float2062Output_2652);

ProductNode_Float2063: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2063weight,ProductNode_Float4Output_5,ProductNode_Float2063Output_2653);

ProductNode_Float2064: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2064weight,ProductNode_Float5Output_6,ProductNode_Float2064Output_2654);

ProductNode_Float2065: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2065weight,vb3,ProductNode_Float2065Output_2655);

ProductNode_Float2066: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2066weight,ProductNode_Float7Output_8,ProductNode_Float2066Output_2656);

ProductNode_Float2067: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2067weight,ProductNode_Float8Output_9,ProductNode_Float2067Output_2657);

SumNode_Float590: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float61Output_73,ProductNode_Float58Output_70,SumNode_Float590Output_2658);

ProductNode_Float2068: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float12Output_74,ProductNode_Float55Output_67,ProductNode_Float2068Output_2659);

ProductNode_Float2069: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2069weight,ProductNode_Float62Output_75,ProductNode_Float2069Output_2660);

ProductNode_Float2070: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2070weight,v8,ProductNode_Float2070Output_2661);

ProductNode_Float2071: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2071weight,vb8,ProductNode_Float2071Output_2662);

SumNode_Float591: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float65Output_78,ProductNode_Float64Output_77,SumNode_Float591Output_2663);

ProductNode_Float2072: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb7,SumNode_Float13Output_79,ProductNode_Float2072Output_2664);

ProductNode_Float2073: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2073weight,v3,ProductNode_Float2073Output_2665);

ProductNode_Float2074: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2074weight,ProductNode_Float4Output_5,ProductNode_Float2074Output_2666);

ProductNode_Float2075: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2075weight,ProductNode_Float16Output_19,ProductNode_Float2075Output_2667);

ProductNode_Float2076: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2076weight,vb3,ProductNode_Float2076Output_2668);

ProductNode_Float2077: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2077weight,ProductNode_Float7Output_8,ProductNode_Float2077Output_2669);

ProductNode_Float2078: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2078weight,ProductNode_Float19Output_22,ProductNode_Float2078Output_2670);

SumNode_Float592: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float72Output_86,ProductNode_Float69Output_83,SumNode_Float592Output_2671);

ProductNode_Float2079: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float14Output_87,ProductNode_Float66Output_80,ProductNode_Float2079Output_2672);

ProductNode_Float2080: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2080weight,ProductNode_Float73Output_88,ProductNode_Float2080Output_2673);

SumNode_Float593: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float647Output_827,ProductNode_Float636Output_814,SumNode_Float593Output_2674);

ProductNode_Float2081: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float180Output_828,ProductNode_Float0Output_0,ProductNode_Float2081Output_2675);

ProductNode_Float2082: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2082weight,ProductNode_Float648Output_829,ProductNode_Float2082Output_2676);

ProductNode_Float2083: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2083weight,vb4,ProductNode_Float2083Output_2677);

ProductNode_Float2084: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2084weight,v8,ProductNode_Float2084Output_2678);

ProductNode_Float2085: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2085weight,vb8,ProductNode_Float2085Output_2679);

SumNode_Float594: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float79Output_95,ProductNode_Float78Output_94,SumNode_Float594Output_2680);

ProductNode_Float2086: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v7,SumNode_Float16Output_96,ProductNode_Float2086Output_2681);

ProductNode_Float2087: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2087weight,v3,ProductNode_Float2087Output_2682);

ProductNode_Float2088: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2088weight,ProductNode_Float29Output_35,ProductNode_Float2088Output_2683);

ProductNode_Float2089: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2089weight,ProductNode_Float30Output_36,ProductNode_Float2089Output_2684);

ProductNode_Float2090: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2090weight,vb3,ProductNode_Float2090Output_2685);

ProductNode_Float2091: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2091weight,ProductNode_Float32Output_38,ProductNode_Float2091Output_2686);

ProductNode_Float2092: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2092weight,ProductNode_Float33Output_39,ProductNode_Float2092Output_2687);

SumNode_Float595: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float86Output_103,ProductNode_Float83Output_100,SumNode_Float595Output_2688);

ProductNode_Float2093: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float17Output_104,ProductNode_Float80Output_97,ProductNode_Float2093Output_2689);

ProductNode_Float2094: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2094weight,ProductNode_Float87Output_105,ProductNode_Float2094Output_2690);

ProductNode_Float2095: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2095weight,v8,ProductNode_Float2095Output_2691);

ProductNode_Float2096: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2096weight,vb8,ProductNode_Float2096Output_2692);

SumNode_Float596: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float90Output_108,ProductNode_Float89Output_107,SumNode_Float596Output_2693);

ProductNode_Float2097: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb7,SumNode_Float18Output_109,ProductNode_Float2097Output_2694);

ProductNode_Float2098: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2098weight,v3,ProductNode_Float2098Output_2695);

ProductNode_Float2099: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2099weight,ProductNode_Float29Output_35,ProductNode_Float2099Output_2696);

ProductNode_Float2100: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2100weight,ProductNode_Float41Output_49,ProductNode_Float2100Output_2697);

ProductNode_Float2101: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2101weight,vb3,ProductNode_Float2101Output_2698);

ProductNode_Float2102: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2102weight,ProductNode_Float32Output_38,ProductNode_Float2102Output_2699);

ProductNode_Float2103: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2103weight,ProductNode_Float44Output_52,ProductNode_Float2103Output_2700);

SumNode_Float597: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float97Output_116,ProductNode_Float94Output_113,SumNode_Float597Output_2701);

ProductNode_Float2104: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float19Output_117,ProductNode_Float91Output_110,ProductNode_Float2104Output_2702);

ProductNode_Float2105: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2105weight,ProductNode_Float98Output_118,ProductNode_Float2105Output_2703);

SumNode_Float598: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float672Output_857,ProductNode_Float661Output_844,SumNode_Float598Output_2704);

ProductNode_Float2106: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float185Output_858,ProductNode_Float25Output_30,ProductNode_Float2106Output_2705);

ProductNode_Float2107: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2107weight,ProductNode_Float673Output_859,ProductNode_Float2107Output_2706);

SumNode_Float599: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float960Output_1228,ProductNode_Float935Output_1198,SumNode_Float599Output_2707);

ProductNode_Float2108: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb5,SumNode_Float268Output_1229,ProductNode_Float2108Output_2708);

ProductNode_Float2109: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2109weight,ProductNode_Float961Output_1230,ProductNode_Float2109Output_2709);

SumNode_Float600: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2109Output_2709,ProductNode_Float2057Output_2646,SumNode_Float600Output_2710);

ProductNode_Float2110: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb16,SumNode_Float600Output_2710,ProductNode_Float2110Output_2711);

ProductNode_Float2111: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2111weight,v11,ProductNode_Float2111Output_2712);

ProductNode_Float2112: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2112weight,vb11,ProductNode_Float2112Output_2713);

SumNode_Float601: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float679Output_867,ProductNode_Float678Output_866,SumNode_Float601Output_2714);

ProductNode_Float2113: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v12,SumNode_Float188Output_868,ProductNode_Float2113Output_2715);

ProductNode_Float2114: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2114weight,ProductNode_Float680Output_869,ProductNode_Float2114Output_2716);

ProductNode_Float2115: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2115weight,v2,ProductNode_Float2115Output_2717);

ProductNode_Float2116: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2116weight,vb2,ProductNode_Float2116Output_2718);

SumNode_Float602: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float110Output_134,ProductNode_Float109Output_133,SumNode_Float602Output_2719);

ProductNode_Float2117: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float24Output_135,ProductNode_Float681Output_870,ProductNode_Float2117Output_2720);

ProductNode_Float2118: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2118weight,v11,ProductNode_Float2118Output_2721);

ProductNode_Float2119: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2119weight,vb11,ProductNode_Float2119Output_2722);

SumNode_Float603: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float686Output_876,ProductNode_Float685Output_875,SumNode_Float603Output_2723);

ProductNode_Float2120: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb12,SumNode_Float190Output_877,ProductNode_Float2120Output_2724);

ProductNode_Float2121: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2121weight,ProductNode_Float687Output_878,ProductNode_Float2121Output_2725);

ProductNode_Float2122: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2122weight,v2,ProductNode_Float2122Output_2726);

ProductNode_Float2123: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2123weight,vb2,ProductNode_Float2123Output_2727);

SumNode_Float604: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float117Output_143,ProductNode_Float116Output_142,SumNode_Float604Output_2728);

ProductNode_Float2124: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float26Output_144,ProductNode_Float688Output_879,ProductNode_Float2124Output_2729);

SumNode_Float605: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float691Output_883,ProductNode_Float684Output_874,SumNode_Float605Output_2730);

ProductNode_Float2125: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v13,SumNode_Float192Output_884,ProductNode_Float2125Output_2731);

ProductNode_Float2126: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2126weight,ProductNode_Float692Output_885,ProductNode_Float2126Output_2732);

ProductNode_Float2127: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2127weight,v11,ProductNode_Float2127Output_2733);

ProductNode_Float2128: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2128weight,vb11,ProductNode_Float2128Output_2734);

SumNode_Float606: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float695Output_888,ProductNode_Float694Output_887,SumNode_Float606Output_2735);

ProductNode_Float2129: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v12,SumNode_Float193Output_889,ProductNode_Float2129Output_2736);

ProductNode_Float2130: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2130weight,ProductNode_Float696Output_890,ProductNode_Float2130Output_2737);

ProductNode_Float2131: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2131weight,v2,ProductNode_Float2131Output_2738);

ProductNode_Float2132: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2132weight,vb2,ProductNode_Float2132Output_2739);

SumNode_Float607: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float126Output_155,ProductNode_Float125Output_154,SumNode_Float607Output_2740);

ProductNode_Float2133: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float29Output_156,ProductNode_Float697Output_891,ProductNode_Float2133Output_2741);

ProductNode_Float2134: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2134weight,v11,ProductNode_Float2134Output_2742);

ProductNode_Float2135: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2135weight,vb11,ProductNode_Float2135Output_2743);

SumNode_Float608: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float702Output_897,ProductNode_Float701Output_896,SumNode_Float608Output_2744);

ProductNode_Float2136: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb12,SumNode_Float195Output_898,ProductNode_Float2136Output_2745);

ProductNode_Float2137: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2137weight,ProductNode_Float703Output_899,ProductNode_Float2137Output_2746);

ProductNode_Float2138: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2138weight,v2,ProductNode_Float2138Output_2747);

ProductNode_Float2139: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2139weight,vb2,ProductNode_Float2139Output_2748);

SumNode_Float609: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float133Output_164,ProductNode_Float132Output_163,SumNode_Float609Output_2749);

ProductNode_Float2140: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float31Output_165,ProductNode_Float704Output_900,ProductNode_Float2140Output_2750);

SumNode_Float610: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float707Output_904,ProductNode_Float700Output_895,SumNode_Float610Output_2751);

ProductNode_Float2141: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb13,SumNode_Float197Output_905,ProductNode_Float2141Output_2752);

ProductNode_Float2142: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2142weight,ProductNode_Float708Output_906,ProductNode_Float2142Output_2753);

SumNode_Float611: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float709Output_907,ProductNode_Float693Output_886,SumNode_Float611Output_2754);

ProductNode_Float2143: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v10,SumNode_Float198Output_908,ProductNode_Float2143Output_2755);

ProductNode_Float2144: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2144weight,v1,ProductNode_Float2144Output_2756);

ProductNode_Float2145: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2145weight,vb1,ProductNode_Float2145Output_2757);

SumNode_Float612: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1286Output_1651,ProductNode_Float1285Output_1650,SumNode_Float612Output_2758);

ProductNode_Float2146: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v9,SumNode_Float365Output_1652,ProductNode_Float2146Output_2759);

ProductNode_Float2147: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2147weight,ProductNode_Float1287Output_1653,ProductNode_Float2147Output_2760);

ProductNode_Float2148: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2148weight,ProductNode_Float1288Output_1654,ProductNode_Float2148Output_2761);

ProductNode_Float2149: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2149weight,v1,ProductNode_Float2149Output_2762);

ProductNode_Float2150: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2150weight,vb1,ProductNode_Float2150Output_2763);

SumNode_Float613: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1291Output_1657,ProductNode_Float1290Output_1656,SumNode_Float613Output_2764);

ProductNode_Float2151: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb9,SumNode_Float366Output_1658,ProductNode_Float2151Output_2765);

ProductNode_Float2152: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2152weight,ProductNode_Float1292Output_1659,ProductNode_Float2152Output_2766);

ProductNode_Float2153: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2153weight,ProductNode_Float1293Output_1660,ProductNode_Float2153Output_2767);

SumNode_Float614: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1294Output_1661,ProductNode_Float1289Output_1655,SumNode_Float614Output_2768);

ProductNode_Float2154: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float367Output_1662,ProductNode_Float710Output_909,ProductNode_Float2154Output_2769);

ProductNode_Float2155: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2155weight,v11,ProductNode_Float2155Output_2770);

ProductNode_Float2156: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2156weight,vb11,ProductNode_Float2156Output_2771);

SumNode_Float615: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float679Output_867,ProductNode_Float678Output_866,SumNode_Float615Output_2772);

ProductNode_Float2157: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v12,SumNode_Float188Output_868,ProductNode_Float2157Output_2773);

ProductNode_Float2158: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2158weight,ProductNode_Float680Output_869,ProductNode_Float2158Output_2774);

ProductNode_Float2159: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2159weight,v2,ProductNode_Float2159Output_2775);

ProductNode_Float2160: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2160weight,vb2,ProductNode_Float2160Output_2776);

SumNode_Float616: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float110Output_134,ProductNode_Float109Output_133,SumNode_Float616Output_2777);

ProductNode_Float2161: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float24Output_135,ProductNode_Float681Output_870,ProductNode_Float2161Output_2778);

ProductNode_Float2162: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2162weight,v11,ProductNode_Float2162Output_2779);

ProductNode_Float2163: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2163weight,vb11,ProductNode_Float2163Output_2780);

SumNode_Float617: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float686Output_876,ProductNode_Float685Output_875,SumNode_Float617Output_2781);

ProductNode_Float2164: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb12,SumNode_Float190Output_877,ProductNode_Float2164Output_2782);

ProductNode_Float2165: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2165weight,ProductNode_Float687Output_878,ProductNode_Float2165Output_2783);

ProductNode_Float2166: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2166weight,v2,ProductNode_Float2166Output_2784);

ProductNode_Float2167: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2167weight,vb2,ProductNode_Float2167Output_2785);

SumNode_Float618: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float117Output_143,ProductNode_Float116Output_142,SumNode_Float618Output_2786);

ProductNode_Float2168: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float26Output_144,ProductNode_Float688Output_879,ProductNode_Float2168Output_2787);

SumNode_Float619: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float691Output_883,ProductNode_Float684Output_874,SumNode_Float619Output_2788);

ProductNode_Float2169: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v13,SumNode_Float192Output_884,ProductNode_Float2169Output_2789);

ProductNode_Float2170: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2170weight,ProductNode_Float692Output_885,ProductNode_Float2170Output_2790);

ProductNode_Float2171: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2171weight,v11,ProductNode_Float2171Output_2791);

ProductNode_Float2172: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2172weight,vb11,ProductNode_Float2172Output_2792);

SumNode_Float620: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float695Output_888,ProductNode_Float694Output_887,SumNode_Float620Output_2793);

ProductNode_Float2173: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v12,SumNode_Float193Output_889,ProductNode_Float2173Output_2794);

ProductNode_Float2174: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2174weight,ProductNode_Float696Output_890,ProductNode_Float2174Output_2795);

ProductNode_Float2175: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2175weight,v2,ProductNode_Float2175Output_2796);

ProductNode_Float2176: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2176weight,vb2,ProductNode_Float2176Output_2797);

SumNode_Float621: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float126Output_155,ProductNode_Float125Output_154,SumNode_Float621Output_2798);

ProductNode_Float2177: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float29Output_156,ProductNode_Float697Output_891,ProductNode_Float2177Output_2799);

ProductNode_Float2178: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2178weight,v11,ProductNode_Float2178Output_2800);

ProductNode_Float2179: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2179weight,vb11,ProductNode_Float2179Output_2801);

SumNode_Float622: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float702Output_897,ProductNode_Float701Output_896,SumNode_Float622Output_2802);

ProductNode_Float2180: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb12,SumNode_Float195Output_898,ProductNode_Float2180Output_2803);

ProductNode_Float2181: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2181weight,ProductNode_Float703Output_899,ProductNode_Float2181Output_2804);

ProductNode_Float2182: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2182weight,v2,ProductNode_Float2182Output_2805);

ProductNode_Float2183: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2183weight,vb2,ProductNode_Float2183Output_2806);

SumNode_Float623: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float133Output_164,ProductNode_Float132Output_163,SumNode_Float623Output_2807);

ProductNode_Float2184: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float31Output_165,ProductNode_Float704Output_900,ProductNode_Float2184Output_2808);

SumNode_Float624: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float707Output_904,ProductNode_Float700Output_895,SumNode_Float624Output_2809);

ProductNode_Float2185: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb13,SumNode_Float197Output_905,ProductNode_Float2185Output_2810);

ProductNode_Float2186: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2186weight,ProductNode_Float708Output_906,ProductNode_Float2186Output_2811);

SumNode_Float625: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float753Output_965,ProductNode_Float737Output_944,SumNode_Float625Output_2812);

ProductNode_Float2187: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb10,SumNode_Float212Output_966,ProductNode_Float2187Output_2813);

ProductNode_Float2188: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2188weight,v1,ProductNode_Float2188Output_2814);

ProductNode_Float2189: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2189weight,vb1,ProductNode_Float2189Output_2815);

SumNode_Float626: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1330Output_1709,ProductNode_Float1329Output_1708,SumNode_Float626Output_2816);

ProductNode_Float2190: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v9,SumNode_Float379Output_1710,ProductNode_Float2190Output_2817);

ProductNode_Float2191: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2191weight,ProductNode_Float1331Output_1711,ProductNode_Float2191Output_2818);

ProductNode_Float2192: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2192weight,ProductNode_Float1332Output_1712,ProductNode_Float2192Output_2819);

ProductNode_Float2193: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2193weight,v1,ProductNode_Float2193Output_2820);

ProductNode_Float2194: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2194weight,vb1,ProductNode_Float2194Output_2821);

SumNode_Float627: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1335Output_1715,ProductNode_Float1334Output_1714,SumNode_Float627Output_2822);

ProductNode_Float2195: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb9,SumNode_Float380Output_1716,ProductNode_Float2195Output_2823);

ProductNode_Float2196: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2196weight,ProductNode_Float1336Output_1717,ProductNode_Float2196Output_2824);

ProductNode_Float2197: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2197weight,ProductNode_Float1337Output_1718,ProductNode_Float2197Output_2825);

SumNode_Float628: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1338Output_1719,ProductNode_Float1333Output_1713,SumNode_Float628Output_2826);

ProductNode_Float2198: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float381Output_1720,ProductNode_Float754Output_967,ProductNode_Float2198Output_2827);

SumNode_Float629: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1912Output_2459,ProductNode_Float1868Output_2401,SumNode_Float629Output_2828);

ProductNode_Float2199: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v15,SumNode_Float547Output_2460,ProductNode_Float2199Output_2829);

ProductNode_Float2200: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2200weight,ProductNode_Float1913Output_2461,ProductNode_Float2200Output_2830);

ProductNode_Float2201: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2201weight,v11,ProductNode_Float2201Output_2831);

ProductNode_Float2202: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2202weight,vb11,ProductNode_Float2202Output_2832);

SumNode_Float630: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float679Output_867,ProductNode_Float678Output_866,SumNode_Float630Output_2833);

ProductNode_Float2203: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v12,SumNode_Float188Output_868,ProductNode_Float2203Output_2834);

ProductNode_Float2204: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2204weight,ProductNode_Float680Output_869,ProductNode_Float2204Output_2835);

ProductNode_Float2205: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2205weight,v2,ProductNode_Float2205Output_2836);

ProductNode_Float2206: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2206weight,vb2,ProductNode_Float2206Output_2837);

SumNode_Float631: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float200Output_253,ProductNode_Float199Output_252,SumNode_Float631Output_2838);

ProductNode_Float2207: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float53Output_254,ProductNode_Float681Output_870,ProductNode_Float2207Output_2839);

ProductNode_Float2208: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2208weight,v11,ProductNode_Float2208Output_2840);

ProductNode_Float2209: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2209weight,vb11,ProductNode_Float2209Output_2841);

SumNode_Float632: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float686Output_876,ProductNode_Float685Output_875,SumNode_Float632Output_2842);

ProductNode_Float2210: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb12,SumNode_Float190Output_877,ProductNode_Float2210Output_2843);

ProductNode_Float2211: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2211weight,ProductNode_Float687Output_878,ProductNode_Float2211Output_2844);

ProductNode_Float2212: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2212weight,v2,ProductNode_Float2212Output_2845);

ProductNode_Float2213: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2213weight,vb2,ProductNode_Float2213Output_2846);

SumNode_Float633: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float207Output_262,ProductNode_Float206Output_261,SumNode_Float633Output_2847);

ProductNode_Float2214: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float55Output_263,ProductNode_Float688Output_879,ProductNode_Float2214Output_2848);

SumNode_Float634: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float781Output_1002,ProductNode_Float774Output_993,SumNode_Float634Output_2849);

ProductNode_Float2215: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v13,SumNode_Float221Output_1003,ProductNode_Float2215Output_2850);

ProductNode_Float2216: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2216weight,ProductNode_Float782Output_1004,ProductNode_Float2216Output_2851);

ProductNode_Float2217: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2217weight,v11,ProductNode_Float2217Output_2852);

ProductNode_Float2218: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2218weight,vb11,ProductNode_Float2218Output_2853);

SumNode_Float635: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float695Output_888,ProductNode_Float694Output_887,SumNode_Float635Output_2854);

ProductNode_Float2219: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v12,SumNode_Float193Output_889,ProductNode_Float2219Output_2855);

ProductNode_Float2220: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2220weight,ProductNode_Float696Output_890,ProductNode_Float2220Output_2856);

ProductNode_Float2221: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2221weight,v2,ProductNode_Float2221Output_2857);

ProductNode_Float2222: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2222weight,vb2,ProductNode_Float2222Output_2858);

SumNode_Float636: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float216Output_274,ProductNode_Float215Output_273,SumNode_Float636Output_2859);

ProductNode_Float2223: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float58Output_275,ProductNode_Float697Output_891,ProductNode_Float2223Output_2860);

ProductNode_Float2224: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2224weight,v11,ProductNode_Float2224Output_2861);

ProductNode_Float2225: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2225weight,vb11,ProductNode_Float2225Output_2862);

SumNode_Float637: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float702Output_897,ProductNode_Float701Output_896,SumNode_Float637Output_2863);

ProductNode_Float2226: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb12,SumNode_Float195Output_898,ProductNode_Float2226Output_2864);

ProductNode_Float2227: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2227weight,ProductNode_Float703Output_899,ProductNode_Float2227Output_2865);

ProductNode_Float2228: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2228weight,v2,ProductNode_Float2228Output_2866);

ProductNode_Float2229: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2229weight,vb2,ProductNode_Float2229Output_2867);

SumNode_Float638: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float223Output_283,ProductNode_Float222Output_282,SumNode_Float638Output_2868);

ProductNode_Float2230: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float60Output_284,ProductNode_Float704Output_900,ProductNode_Float2230Output_2869);

SumNode_Float639: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float797Output_1023,ProductNode_Float790Output_1014,SumNode_Float639Output_2870);

ProductNode_Float2231: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb13,SumNode_Float226Output_1024,ProductNode_Float2231Output_2871);

ProductNode_Float2232: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2232weight,ProductNode_Float798Output_1025,ProductNode_Float2232Output_2872);

SumNode_Float640: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float799Output_1026,ProductNode_Float783Output_1005,SumNode_Float640Output_2873);

ProductNode_Float2233: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v10,SumNode_Float227Output_1027,ProductNode_Float2233Output_2874);

ProductNode_Float2234: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2234weight,v1,ProductNode_Float2234Output_2875);

ProductNode_Float2235: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2235weight,vb1,ProductNode_Float2235Output_2876);

SumNode_Float641: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1286Output_1651,ProductNode_Float1285Output_1650,SumNode_Float641Output_2877);

ProductNode_Float2236: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v9,SumNode_Float365Output_1652,ProductNode_Float2236Output_2878);

ProductNode_Float2237: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2237weight,ProductNode_Float1287Output_1653,ProductNode_Float2237Output_2879);

ProductNode_Float2238: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2238weight,ProductNode_Float1378Output_1773,ProductNode_Float2238Output_2880);

ProductNode_Float2239: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2239weight,v1,ProductNode_Float2239Output_2881);

ProductNode_Float2240: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2240weight,vb1,ProductNode_Float2240Output_2882);

SumNode_Float642: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1291Output_1657,ProductNode_Float1290Output_1656,SumNode_Float642Output_2883);

ProductNode_Float2241: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb9,SumNode_Float366Output_1658,ProductNode_Float2241Output_2884);

ProductNode_Float2242: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2242weight,ProductNode_Float1292Output_1659,ProductNode_Float2242Output_2885);

ProductNode_Float2243: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2243weight,ProductNode_Float1383Output_1779,ProductNode_Float2243Output_2886);

SumNode_Float643: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1384Output_1780,ProductNode_Float1379Output_1774,SumNode_Float643Output_2887);

ProductNode_Float2244: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float396Output_1781,ProductNode_Float800Output_1028,ProductNode_Float2244Output_2888);

ProductNode_Float2245: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2245weight,v11,ProductNode_Float2245Output_2889);

ProductNode_Float2246: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2246weight,vb11,ProductNode_Float2246Output_2890);

SumNode_Float644: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float679Output_867,ProductNode_Float678Output_866,SumNode_Float644Output_2891);

ProductNode_Float2247: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v12,SumNode_Float188Output_868,ProductNode_Float2247Output_2892);

ProductNode_Float2248: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2248weight,ProductNode_Float680Output_869,ProductNode_Float2248Output_2893);

ProductNode_Float2249: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2249weight,v2,ProductNode_Float2249Output_2894);

ProductNode_Float2250: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2250weight,vb2,ProductNode_Float2250Output_2895);

SumNode_Float645: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float200Output_253,ProductNode_Float199Output_252,SumNode_Float645Output_2896);

ProductNode_Float2251: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float53Output_254,ProductNode_Float681Output_870,ProductNode_Float2251Output_2897);

ProductNode_Float2252: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2252weight,v11,ProductNode_Float2252Output_2898);

ProductNode_Float2253: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2253weight,vb11,ProductNode_Float2253Output_2899);

SumNode_Float646: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float686Output_876,ProductNode_Float685Output_875,SumNode_Float646Output_2900);

ProductNode_Float2254: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb12,SumNode_Float190Output_877,ProductNode_Float2254Output_2901);

ProductNode_Float2255: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2255weight,ProductNode_Float687Output_878,ProductNode_Float2255Output_2902);

ProductNode_Float2256: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2256weight,v2,ProductNode_Float2256Output_2903);

ProductNode_Float2257: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2257weight,vb2,ProductNode_Float2257Output_2904);

SumNode_Float647: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float207Output_262,ProductNode_Float206Output_261,SumNode_Float647Output_2905);

ProductNode_Float2258: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float55Output_263,ProductNode_Float688Output_879,ProductNode_Float2258Output_2906);

SumNode_Float648: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float781Output_1002,ProductNode_Float774Output_993,SumNode_Float648Output_2907);

ProductNode_Float2259: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v13,SumNode_Float221Output_1003,ProductNode_Float2259Output_2908);

ProductNode_Float2260: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2260weight,ProductNode_Float782Output_1004,ProductNode_Float2260Output_2909);

ProductNode_Float2261: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2261weight,v11,ProductNode_Float2261Output_2910);

ProductNode_Float2262: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2262weight,vb11,ProductNode_Float2262Output_2911);

SumNode_Float649: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float695Output_888,ProductNode_Float694Output_887,SumNode_Float649Output_2912);

ProductNode_Float2263: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v12,SumNode_Float193Output_889,ProductNode_Float2263Output_2913);

ProductNode_Float2264: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2264weight,ProductNode_Float696Output_890,ProductNode_Float2264Output_2914);

ProductNode_Float2265: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2265weight,v2,ProductNode_Float2265Output_2915);

ProductNode_Float2266: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2266weight,vb2,ProductNode_Float2266Output_2916);

SumNode_Float650: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float216Output_274,ProductNode_Float215Output_273,SumNode_Float650Output_2917);

ProductNode_Float2267: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float58Output_275,ProductNode_Float697Output_891,ProductNode_Float2267Output_2918);

ProductNode_Float2268: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2268weight,v11,ProductNode_Float2268Output_2919);

ProductNode_Float2269: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2269weight,vb11,ProductNode_Float2269Output_2920);

SumNode_Float651: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float702Output_897,ProductNode_Float701Output_896,SumNode_Float651Output_2921);

ProductNode_Float2270: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb12,SumNode_Float195Output_898,ProductNode_Float2270Output_2922);

ProductNode_Float2271: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2271weight,ProductNode_Float703Output_899,ProductNode_Float2271Output_2923);

ProductNode_Float2272: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2272weight,v2,ProductNode_Float2272Output_2924);

ProductNode_Float2273: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2273weight,vb2,ProductNode_Float2273Output_2925);

SumNode_Float652: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float223Output_283,ProductNode_Float222Output_282,SumNode_Float652Output_2926);

ProductNode_Float2274: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float60Output_284,ProductNode_Float704Output_900,ProductNode_Float2274Output_2927);

SumNode_Float653: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float797Output_1023,ProductNode_Float790Output_1014,SumNode_Float653Output_2928);

ProductNode_Float2275: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb13,SumNode_Float226Output_1024,ProductNode_Float2275Output_2929);

ProductNode_Float2276: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2276weight,ProductNode_Float798Output_1025,ProductNode_Float2276Output_2930);

SumNode_Float654: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float843Output_1084,ProductNode_Float827Output_1063,SumNode_Float654Output_2931);

ProductNode_Float2277: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb10,SumNode_Float241Output_1085,ProductNode_Float2277Output_2932);

ProductNode_Float2278: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2278weight,v1,ProductNode_Float2278Output_2933);

ProductNode_Float2279: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2279weight,vb1,ProductNode_Float2279Output_2934);

SumNode_Float655: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1330Output_1709,ProductNode_Float1329Output_1708,SumNode_Float655Output_2935);

ProductNode_Float2280: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(v9,SumNode_Float379Output_1710,ProductNode_Float2280Output_2936);

ProductNode_Float2281: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2281weight,ProductNode_Float1331Output_1711,ProductNode_Float2281Output_2937);

ProductNode_Float2282: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2282weight,ProductNode_Float1422Output_1831,ProductNode_Float2282Output_2938);

ProductNode_Float2283: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2283weight,v1,ProductNode_Float2283Output_2939);

ProductNode_Float2284: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2284weight,vb1,ProductNode_Float2284Output_2940);

SumNode_Float656: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1335Output_1715,ProductNode_Float1334Output_1714,SumNode_Float656Output_2941);

ProductNode_Float2285: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb9,SumNode_Float380Output_1716,ProductNode_Float2285Output_2942);

ProductNode_Float2286: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2286weight,ProductNode_Float1336Output_1717,ProductNode_Float2286Output_2943);

ProductNode_Float2287: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2287weight,ProductNode_Float1427Output_1837,ProductNode_Float2287Output_2944);

SumNode_Float657: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float1428Output_1838,ProductNode_Float1423Output_1832,SumNode_Float657Output_2945);

ProductNode_Float2288: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float410Output_1839,ProductNode_Float844Output_1086,ProductNode_Float2288Output_2946);

SumNode_Float658: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2002Output_2578,ProductNode_Float1958Output_2520,SumNode_Float658Output_2947);

ProductNode_Float2289: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb15,SumNode_Float576Output_2579,ProductNode_Float2289Output_2948);

ProductNode_Float2290: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2290weight,ProductNode_Float2003Output_2580,ProductNode_Float2290Output_2949);

SumNode_Float659: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2290Output_2949,ProductNode_Float2200Output_2830,SumNode_Float659Output_2950);

ProductNode_Float2291: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(SumNode_Float659Output_2950,ProductNode_Float2110Output_2711,ProductNode_Float2291Output_2951);

SumNode_Float660: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2291Output_2951,ProductNode_Float2005Output_2583,SumNode_Float660Output_2952);

ProductNode_Float2292: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb6,SumNode_Float660Output_2952,ProductNode_Float2292Output_2953);

SumNode_Float661: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2292Output_2953,ProductNode_Float1719Output_2215,SumNode_Float661Output_2954);

ProductNode_Float2293: entity work.ProductNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(vb14,SumNode_Float661Output_2954,ProductNode_Float2293Output_2955);

SumNode_Float662: entity work.SumNode_Float(rtl)
generic map(mantissaBits,exponentBits)
port map(ProductNode_Float2293Output_2955,ProductNode_Float1146Output_1477,SumNode_Float662Output_2956);

vout <= SumNode_Float662Output_2956;
 
end architecture;

--------------------------------------------------------------------------------
--                    SmallMultTableP3x3r6XuYu_comb_uid33
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2007-2012)
--------------------------------------------------------------------------------
library ieee; 
use ieee.std_logic_1164.all;
library work;
entity SmallMultTableP3x3r6XuYu_comb_uid33 is
   port ( X : in  std_logic_vector(5 downto 0);
          Y : out  std_logic_vector(5 downto 0)   );
end entity;

architecture arch of SmallMultTableP3x3r6XuYu_comb_uid33 is
signal TableOut :  std_logic_vector(5 downto 0);
begin
  with X select TableOut <= 
   "000000" when "000000",
   "000000" when "000001",
   "000000" when "000010",
   "000000" when "000011",
   "000000" when "000100",
   "000000" when "000101",
   "000000" when "000110",
   "000000" when "000111",
   "000000" when "001000",
   "000001" when "001001",
   "000010" when "001010",
   "000011" when "001011",
   "000100" when "001100",
   "000101" when "001101",
   "000110" when "001110",
   "000111" when "001111",
   "000000" when "010000",
   "000010" when "010001",
   "000100" when "010010",
   "000110" when "010011",
   "001000" when "010100",
   "001010" when "010101",
   "001100" when "010110",
   "001110" when "010111",
   "000000" when "011000",
   "000011" when "011001",
   "000110" when "011010",
   "001001" when "011011",
   "001100" when "011100",
   "001111" when "011101",
   "010010" when "011110",
   "010101" when "011111",
   "000000" when "100000",
   "000100" when "100001",
   "001000" when "100010",
   "001100" when "100011",
   "010000" when "100100",
   "010100" when "100101",
   "011000" when "100110",
   "011100" when "100111",
   "000000" when "101000",
   "000101" when "101001",
   "001010" when "101010",
   "001111" when "101011",
   "010100" when "101100",
   "011001" when "101101",
   "011110" when "101110",
   "100011" when "101111",
   "000000" when "110000",
   "000110" when "110001",
   "001100" when "110010",
   "010010" when "110011",
   "011000" when "110100",
   "011110" when "110101",
   "100100" when "110110",
   "101010" when "110111",
   "000000" when "111000",
   "000111" when "111001",
   "001110" when "111010",
   "010101" when "111011",
   "011100" when "111100",
   "100011" when "111101",
   "101010" when "111110",
   "110001" when "111111",
   "------" when others;
    Y <= TableOut;
end architecture;

--------------------------------------------------------------------------------
--                    SmallMultTableP3x3r6XuYu_comb_uid68
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2007-2012)
--------------------------------------------------------------------------------
library ieee; 
use ieee.std_logic_1164.all;
library work;
entity SmallMultTableP3x3r6XuYu_comb_uid68 is
   port ( X : in  std_logic_vector(5 downto 0);
          Y : out  std_logic_vector(5 downto 0)   );
end entity;

architecture arch of SmallMultTableP3x3r6XuYu_comb_uid68 is
signal TableOut :  std_logic_vector(5 downto 0);
begin
  with X select TableOut <= 
   "000000" when "000000",
   "000000" when "000001",
   "000000" when "000010",
   "000000" when "000011",
   "000000" when "000100",
   "000000" when "000101",
   "000000" when "000110",
   "000000" when "000111",
   "000000" when "001000",
   "000001" when "001001",
   "000010" when "001010",
   "000011" when "001011",
   "000100" when "001100",
   "000101" when "001101",
   "000110" when "001110",
   "000111" when "001111",
   "000000" when "010000",
   "000010" when "010001",
   "000100" when "010010",
   "000110" when "010011",
   "001000" when "010100",
   "001010" when "010101",
   "001100" when "010110",
   "001110" when "010111",
   "000000" when "011000",
   "000011" when "011001",
   "000110" when "011010",
   "001001" when "011011",
   "001100" when "011100",
   "001111" when "011101",
   "010010" when "011110",
   "010101" when "011111",
   "000000" when "100000",
   "000100" when "100001",
   "001000" when "100010",
   "001100" when "100011",
   "010000" when "100100",
   "010100" when "100101",
   "011000" when "100110",
   "011100" when "100111",
   "000000" when "101000",
   "000101" when "101001",
   "001010" when "101010",
   "001111" when "101011",
   "010100" when "101100",
   "011001" when "101101",
   "011110" when "101110",
   "100011" when "101111",
   "000000" when "110000",
   "000110" when "110001",
   "001100" when "110010",
   "010010" when "110011",
   "011000" when "110100",
   "011110" when "110101",
   "100100" when "110110",
   "101010" when "110111",
   "000000" when "111000",
   "000111" when "111001",
   "001110" when "111010",
   "010101" when "111011",
   "011100" when "111100",
   "100011" when "111101",
   "101010" when "111110",
   "110001" when "111111",
   "------" when others;
    Y <= TableOut;
end architecture;

--------------------------------------------------------------------------------
--                    SmallMultTableP3x3r6XuYu_comb_uid103
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin (2007-2012)
--------------------------------------------------------------------------------
library ieee; 
use ieee.std_logic_1164.all;
library work;
entity SmallMultTableP3x3r6XuYu_comb_uid103 is
   port ( X : in  std_logic_vector(5 downto 0);
          Y : out  std_logic_vector(5 downto 0)   );
end entity;

architecture arch of SmallMultTableP3x3r6XuYu_comb_uid103 is
signal TableOut :  std_logic_vector(5 downto 0);
begin
  with X select TableOut <= 
   "000000" when "000000",
   "000000" when "000001",
   "000000" when "000010",
   "000000" when "000011",
   "000000" when "000100",
   "000000" when "000101",
   "000000" when "000110",
   "000000" when "000111",
   "000000" when "001000",
   "000001" when "001001",
   "000010" when "001010",
   "000011" when "001011",
   "000100" when "001100",
   "000101" when "001101",
   "000110" when "001110",
   "000111" when "001111",
   "000000" when "010000",
   "000010" when "010001",
   "000100" when "010010",
   "000110" when "010011",
   "001000" when "010100",
   "001010" when "010101",
   "001100" when "010110",
   "001110" when "010111",
   "000000" when "011000",
   "000011" when "011001",
   "000110" when "011010",
   "001001" when "011011",
   "001100" when "011100",
   "001111" when "011101",
   "010010" when "011110",
   "010101" when "011111",
   "000000" when "100000",
   "000100" when "100001",
   "001000" when "100010",
   "001100" when "100011",
   "010000" when "100100",
   "010100" when "100101",
   "011000" when "100110",
   "011100" when "100111",
   "000000" when "101000",
   "000101" when "101001",
   "001010" when "101010",
   "001111" when "101011",
   "010100" when "101100",
   "011001" when "101101",
   "011110" when "101110",
   "100011" when "101111",
   "000000" when "110000",
   "000110" when "110001",
   "001100" when "110010",
   "010010" when "110011",
   "011000" when "110100",
   "011110" when "110101",
   "100100" when "110110",
   "101010" when "110111",
   "000000" when "111000",
   "000111" when "111001",
   "001110" when "111010",
   "010101" when "111011",
   "011100" when "111100",
   "100011" when "111101",
   "101010" when "111110",
   "110001" when "111111",
   "------" when others;
    Y <= TableOut;
end architecture;

--------------------------------------------------------------------------------
--                               Compressor_6_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Popa, Illyes Kinga, 2012
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_6_3 is
   port ( X0 : in  std_logic_vector(5 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_6_3 is
signal X :  std_logic_vector(5 downto 0);
begin
   X <=X0 ;
   with X select R <= 
      "000" when "000000", 
      "001" when "000001", 
      "001" when "000010", 
      "010" when "000011", 
      "001" when "000100", 
      "010" when "000101", 
      "010" when "000110", 
      "011" when "000111", 
      "001" when "001000", 
      "010" when "001001", 
      "010" when "001010", 
      "011" when "001011", 
      "010" when "001100", 
      "011" when "001101", 
      "011" when "001110", 
      "100" when "001111", 
      "001" when "010000", 
      "010" when "010001", 
      "010" when "010010", 
      "011" when "010011", 
      "010" when "010100", 
      "011" when "010101", 
      "011" when "010110", 
      "100" when "010111", 
      "010" when "011000", 
      "011" when "011001", 
      "011" when "011010", 
      "100" when "011011", 
      "011" when "011100", 
      "100" when "011101", 
      "100" when "011110", 
      "101" when "011111", 
      "001" when "100000", 
      "010" when "100001", 
      "010" when "100010", 
      "011" when "100011", 
      "010" when "100100", 
      "011" when "100101", 
      "011" when "100110", 
      "100" when "100111", 
      "010" when "101000", 
      "011" when "101001", 
      "011" when "101010", 
      "100" when "101011", 
      "011" when "101100", 
      "100" when "101101", 
      "100" when "101110", 
      "101" when "101111", 
      "010" when "110000", 
      "011" when "110001", 
      "011" when "110010", 
      "100" when "110011", 
      "011" when "110100", 
      "100" when "110101", 
      "100" when "110110", 
      "101" when "110111", 
      "011" when "111000", 
      "100" when "111001", 
      "100" when "111010", 
      "101" when "111011", 
      "100" when "111100", 
      "101" when "111101", 
      "101" when "111110", 
      "110" when "111111", 
      "---" when others;

end architecture;

--------------------------------------------------------------------------------
--                              Compressor_14_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Popa, Illyes Kinga, 2012
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_14_3 is
   port ( X0 : in  std_logic_vector(3 downto 0);
          X1 : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_14_3 is
signal X :  std_logic_vector(4 downto 0);
begin
   X <=X1 & X0 ;
   with X select R <= 
      "000" when "00000", 
      "001" when "00001", 
      "001" when "00010", 
      "010" when "00011", 
      "001" when "00100", 
      "010" when "00101", 
      "010" when "00110", 
      "011" when "00111", 
      "001" when "01000", 
      "010" when "01001", 
      "010" when "01010", 
      "011" when "01011", 
      "010" when "01100", 
      "011" when "01101", 
      "011" when "01110", 
      "100" when "01111", 
      "010" when "10000", 
      "011" when "10001", 
      "011" when "10010", 
      "100" when "10011", 
      "011" when "10100", 
      "100" when "10101", 
      "100" when "10110", 
      "101" when "10111", 
      "011" when "11000", 
      "100" when "11001", 
      "100" when "11010", 
      "101" when "11011", 
      "100" when "11100", 
      "101" when "11101", 
      "101" when "11110", 
      "110" when "11111", 
      "---" when others;

end architecture;

--------------------------------------------------------------------------------
--                               Compressor_5_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Popa, Illyes Kinga, 2012
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_5_3 is
   port ( X0 : in  std_logic_vector(4 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_5_3 is
signal X :  std_logic_vector(4 downto 0);
begin
   X <=X0 ;
   with X select R <= 
      "000" when "00000", 
      "001" when "00001", 
      "001" when "00010", 
      "010" when "00011", 
      "001" when "00100", 
      "010" when "00101", 
      "010" when "00110", 
      "011" when "00111", 
      "001" when "01000", 
      "010" when "01001", 
      "010" when "01010", 
      "011" when "01011", 
      "010" when "01100", 
      "011" when "01101", 
      "011" when "01110", 
      "100" when "01111", 
      "001" when "10000", 
      "010" when "10001", 
      "010" when "10010", 
      "011" when "10011", 
      "010" when "10100", 
      "011" when "10101", 
      "011" when "10110", 
      "100" when "10111", 
      "010" when "11000", 
      "011" when "11001", 
      "011" when "11010", 
      "100" when "11011", 
      "011" when "11100", 
      "100" when "11101", 
      "100" when "11110", 
      "101" when "11111", 
      "---" when others;

end architecture;

--------------------------------------------------------------------------------
--                               Compressor_4_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Popa, Illyes Kinga, 2012
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_4_3 is
   port ( X0 : in  std_logic_vector(3 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_4_3 is
signal X :  std_logic_vector(3 downto 0);
begin
   X <=X0 ;
   with X select R <= 
      "000" when "0000", 
      "001" when "0001", 
      "001" when "0010", 
      "010" when "0011", 
      "001" when "0100", 
      "010" when "0101", 
      "010" when "0110", 
      "011" when "0111", 
      "001" when "1000", 
      "010" when "1001", 
      "010" when "1010", 
      "011" when "1011", 
      "010" when "1100", 
      "011" when "1101", 
      "011" when "1110", 
      "100" when "1111", 
      "---" when others;

end architecture;

--------------------------------------------------------------------------------
--                              Compressor_23_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Popa, Illyes Kinga, 2012
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_23_3 is
   port ( X0 : in  std_logic_vector(2 downto 0);
          X1 : in  std_logic_vector(1 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_23_3 is
signal X :  std_logic_vector(4 downto 0);
begin
   X <=X1 & X0 ;
   with X select R <= 
      "000" when "00000", 
      "001" when "00001", 
      "001" when "00010", 
      "010" when "00011", 
      "001" when "00100", 
      "010" when "00101", 
      "010" when "00110", 
      "011" when "00111", 
      "010" when "01000", 
      "011" when "01001", 
      "011" when "01010", 
      "100" when "01011", 
      "011" when "01100", 
      "100" when "01101", 
      "100" when "01110", 
      "101" when "01111", 
      "010" when "10000", 
      "011" when "10001", 
      "011" when "10010", 
      "100" when "10011", 
      "011" when "10100", 
      "100" when "10101", 
      "100" when "10110", 
      "101" when "10111", 
      "100" when "11000", 
      "101" when "11001", 
      "101" when "11010", 
      "110" when "11011", 
      "101" when "11100", 
      "110" when "11101", 
      "110" when "11110", 
      "111" when "11111", 
      "---" when others;

end architecture;

--------------------------------------------------------------------------------
--                              Compressor_13_3
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Popa, Illyes Kinga, 2012
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_13_3 is
   port ( X0 : in  std_logic_vector(2 downto 0);
          X1 : in  std_logic_vector(0 downto 0);
          R : out  std_logic_vector(2 downto 0)   );
end entity;

architecture arch of Compressor_13_3 is
signal X :  std_logic_vector(3 downto 0);
begin
   X <=X1 & X0 ;
   with X select R <= 
      "000" when "0000", 
      "001" when "0001", 
      "001" when "0010", 
      "010" when "0011", 
      "001" when "0100", 
      "010" when "0101", 
      "010" when "0110", 
      "011" when "0111", 
      "010" when "1000", 
      "011" when "1001", 
      "011" when "1010", 
      "100" when "1011", 
      "011" when "1100", 
      "100" when "1101", 
      "100" when "1110", 
      "101" when "1111", 
      "---" when others;

end architecture;

--------------------------------------------------------------------------------
--                               Compressor_3_2
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Popa, Illyes Kinga, 2012
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity Compressor_3_2 is
   port ( X0 : in  std_logic_vector(2 downto 0);
          R : out  std_logic_vector(1 downto 0)   );
end entity;

architecture arch of Compressor_3_2 is
signal X :  std_logic_vector(2 downto 0);
begin
   X <=X0 ;
   with X select R <= 
      "00" when "000", 
      "01" when "001", 
      "01" when "010", 
      "10" when "011", 
      "01" when "100", 
      "10" when "101", 
      "10" when "110", 
      "11" when "111", 
      "--" when others;

end architecture;

--------------------------------------------------------------------------------
--                             LZOC_64_comb_uid6
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007)
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LZOC_64_comb_uid6 is
   port ( I : in  std_logic_vector(63 downto 0);
          OZB : in  std_logic;
          O : out  std_logic_vector(6 downto 0)   );
end entity;

architecture arch of LZOC_64_comb_uid6 is
signal sozb :  std_logic;
signal level7 :  std_logic_vector(127 downto 0);
signal digit7 :  std_logic;
signal level6 :  std_logic_vector(63 downto 0);
signal digit6 :  std_logic;
signal level5 :  std_logic_vector(31 downto 0);
signal digit5 :  std_logic;
signal level4 :  std_logic_vector(15 downto 0);
signal digit4 :  std_logic;
signal level3 :  std_logic_vector(7 downto 0);
signal digit3 :  std_logic;
signal level2 :  std_logic_vector(3 downto 0);
signal digit2 :  std_logic;
signal level1 :  std_logic_vector(1 downto 0);
signal digit1 :  std_logic;
begin
   sozb <= OZB;
   level7<= I& (63 downto 0 => not(sozb));
   digit7<= '1' when level7(127 downto 64) = (127 downto 64 => sozb) else '0';
   level6<= level7(63 downto 0) when digit7='1' else level7(127 downto 64);
   digit6<= '1' when level6(63 downto 32) = (63 downto 32 => sozb) else '0';
   level5<= level6(31 downto 0) when digit6='1' else level6(63 downto 32);
   digit5<= '1' when level5(31 downto 16) = (31 downto 16 => sozb) else '0';
   level4<= level5(15 downto 0) when digit5='1' else level5(31 downto 16);
   digit4<= '1' when level4(15 downto 8) = (15 downto 8 => sozb) else '0';
   level3<= level4(7 downto 0) when digit4='1' else level4(15 downto 8);
   digit3<= '1' when level3(7 downto 4) = (7 downto 4 => sozb) else '0';
   level2<= level3(3 downto 0) when digit3='1' else level3(7 downto 4);
   digit2<= '1' when level2(3 downto 2) = (3 downto 2 => sozb) else '0';
   level1<= level2(1 downto 0) when digit2='1' else level2(3 downto 2);
   digit1<= '1' when level1(1 downto 1) = (1 downto 1 => sozb) else '0';
   O <= digit7 & digit6 & digit5 & digit4 & digit3 & digit2 & digit1;
end architecture;

--------------------------------------------------------------------------------
--                    LeftShifter_64_by_max_64_comb_uid10
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2011)
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LeftShifter_64_by_max_64_comb_uid10 is
   port ( X : in  std_logic_vector(63 downto 0);
          S : in  std_logic_vector(6 downto 0);
          R : out  std_logic_vector(127 downto 0)   );
end entity;

architecture arch of LeftShifter_64_by_max_64_comb_uid10 is
signal level0 :  std_logic_vector(63 downto 0);
signal ps :  std_logic_vector(6 downto 0);
signal level1 :  std_logic_vector(64 downto 0);
signal level2 :  std_logic_vector(66 downto 0);
signal level3 :  std_logic_vector(70 downto 0);
signal level4 :  std_logic_vector(78 downto 0);
signal level5 :  std_logic_vector(94 downto 0);
signal level6 :  std_logic_vector(126 downto 0);
signal level7 :  std_logic_vector(190 downto 0);
begin
   level0<= X;
   ps<= S;
   level1<= level0 & (0 downto 0 => '0') when ps(0)= '1' else     (0 downto 0 => '0') & level0;
   level2<= level1 & (1 downto 0 => '0') when ps(1)= '1' else     (1 downto 0 => '0') & level1;
   level3<= level2 & (3 downto 0 => '0') when ps(2)= '1' else     (3 downto 0 => '0') & level2;
   level4<= level3 & (7 downto 0 => '0') when ps(3)= '1' else     (7 downto 0 => '0') & level3;
   level5<= level4 & (15 downto 0 => '0') when ps(4)= '1' else     (15 downto 0 => '0') & level4;
   level6<= level5 & (31 downto 0 => '0') when ps(5)= '1' else     (31 downto 0 => '0') & level5;
   level7<= level6 & (63 downto 0 => '0') when ps(6)= '1' else     (63 downto 0 => '0') & level6;
   R <= level7(127 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                        PositDecoder_65_7_comb_uid4
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Raul Murillo, 2019
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity PositDecoder_65_7_comb_uid4 is
   port ( Input : in  std_logic_vector(64 downto 0);
          Sign : out  std_logic;
          Reg : out  std_logic_vector(7 downto 0);
          Exp : out  std_logic_vector(6 downto 0);
          Frac : out  std_logic_vector(55 downto 0);
          z : out  std_logic;
          inf : out  std_logic   );
end entity;

architecture arch of PositDecoder_65_7_comb_uid4 is
   component LZOC_64_comb_uid6 is
      port ( I : in  std_logic_vector(63 downto 0);
             OZB : in  std_logic;
             O : out  std_logic_vector(6 downto 0)   );
   end component;

   component LeftShifter_64_by_max_64_comb_uid10 is
      port ( X : in  std_logic_vector(63 downto 0);
             S : in  std_logic_vector(6 downto 0);
             R : out  std_logic_vector(127 downto 0)   );
   end component;

signal nzero :  std_logic;
signal my_sign :  std_logic;
signal rep_sign :  std_logic_vector(63 downto 0);
signal twos :  std_logic_vector(63 downto 0);
signal rc :  std_logic;
signal rep_rc :  std_logic_vector(63 downto 0);
signal inv :  std_logic_vector(63 downto 0);
signal zero_var :  std_logic;
signal zc :  std_logic_vector(6 downto 0);
signal zc_sub :  std_logic_vector(6 downto 0);
signal shifted_twos :  std_logic_vector(127 downto 0);
signal tmp :  std_logic_vector(61 downto 0);
begin
-------------------------------- Special Cases --------------------------------
   nzero <= '0' when Input(63 downto 0) = 0 else '1';
   -- 1 if Input is zero
   z <= Input(64) NOR nzero;
   -- 1 if Input is infinity
   inf <= Input(64) AND (NOT nzero);
------------------------------- Extract Sign bit -------------------------------
   my_sign <= Input(64);
   Sign <= my_sign;
--------------------------- 2's Complement of Input ---------------------------
   rep_sign <= (others => my_sign);
   twos <= (rep_sign XOR Input(63 downto 0)) + my_sign;
   rc <= twos(63);
------------------------ Count leading zeros of regime ------------------------
   rep_rc <= (others => rc);
   -- Invert 2's
   inv <= rep_rc XOR twos;
   zero_var <= '0';
   LZOC_Component: LZOC_64_comb_uid6
      port map ( I => inv,
                 O => zc,
                 OZB => zero_var);
----------------------------- Shift out the regime -----------------------------
   zc_sub <= zc - 1;
   LeftShifterComponent: LeftShifter_64_by_max_64_comb_uid10
      port map ( R => shifted_twos,
                 S => zc_sub,
                 X => twos);
   tmp <= shifted_twos(61 downto 0);
------------------------ Extract fraction and exponent ------------------------
   Frac <= nzero & tmp(54 downto 0);
   Exp <= tmp(61 downto 55);
-------------------------------- Select regime --------------------------------
   Reg <= '0' & zc_sub when rc = '1' else NOT('0' & zc) + 1;
end architecture;

--------------------------------------------------------------------------------
--                             LZOC_64_comb_uid18
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Bogdan Pasca (2007)
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LZOC_64_comb_uid18 is
   port ( I : in  std_logic_vector(63 downto 0);
          OZB : in  std_logic;
          O : out  std_logic_vector(6 downto 0)   );
end entity;

architecture arch of LZOC_64_comb_uid18 is
signal sozb :  std_logic;
signal level7 :  std_logic_vector(127 downto 0);
signal digit7 :  std_logic;
signal level6 :  std_logic_vector(63 downto 0);
signal digit6 :  std_logic;
signal level5 :  std_logic_vector(31 downto 0);
signal digit5 :  std_logic;
signal level4 :  std_logic_vector(15 downto 0);
signal digit4 :  std_logic;
signal level3 :  std_logic_vector(7 downto 0);
signal digit3 :  std_logic;
signal level2 :  std_logic_vector(3 downto 0);
signal digit2 :  std_logic;
signal level1 :  std_logic_vector(1 downto 0);
signal digit1 :  std_logic;
begin
   sozb <= OZB;
   level7<= I& (63 downto 0 => not(sozb));
   digit7<= '1' when level7(127 downto 64) = (127 downto 64 => sozb) else '0';
   level6<= level7(63 downto 0) when digit7='1' else level7(127 downto 64);
   digit6<= '1' when level6(63 downto 32) = (63 downto 32 => sozb) else '0';
   level5<= level6(31 downto 0) when digit6='1' else level6(63 downto 32);
   digit5<= '1' when level5(31 downto 16) = (31 downto 16 => sozb) else '0';
   level4<= level5(15 downto 0) when digit5='1' else level5(31 downto 16);
   digit4<= '1' when level4(15 downto 8) = (15 downto 8 => sozb) else '0';
   level3<= level4(7 downto 0) when digit4='1' else level4(15 downto 8);
   digit3<= '1' when level3(7 downto 4) = (7 downto 4 => sozb) else '0';
   level2<= level3(3 downto 0) when digit3='1' else level3(7 downto 4);
   digit2<= '1' when level2(3 downto 2) = (3 downto 2 => sozb) else '0';
   level1<= level2(1 downto 0) when digit2='1' else level2(3 downto 2);
   digit1<= '1' when level1(1 downto 1) = (1 downto 1 => sozb) else '0';
   O <= digit7 & digit6 & digit5 & digit4 & digit3 & digit2 & digit1;
end architecture;

--------------------------------------------------------------------------------
--                    LeftShifter_64_by_max_64_comb_uid22
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2011)
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity LeftShifter_64_by_max_64_comb_uid22 is
   port ( X : in  std_logic_vector(63 downto 0);
          S : in  std_logic_vector(6 downto 0);
          R : out  std_logic_vector(127 downto 0)   );
end entity;

architecture arch of LeftShifter_64_by_max_64_comb_uid22 is
signal level0 :  std_logic_vector(63 downto 0);
signal ps :  std_logic_vector(6 downto 0);
signal level1 :  std_logic_vector(64 downto 0);
signal level2 :  std_logic_vector(66 downto 0);
signal level3 :  std_logic_vector(70 downto 0);
signal level4 :  std_logic_vector(78 downto 0);
signal level5 :  std_logic_vector(94 downto 0);
signal level6 :  std_logic_vector(126 downto 0);
signal level7 :  std_logic_vector(190 downto 0);
begin
   level0<= X;
   ps<= S;
   level1<= level0 & (0 downto 0 => '0') when ps(0)= '1' else     (0 downto 0 => '0') & level0;
   level2<= level1 & (1 downto 0 => '0') when ps(1)= '1' else     (1 downto 0 => '0') & level1;
   level3<= level2 & (3 downto 0 => '0') when ps(2)= '1' else     (3 downto 0 => '0') & level2;
   level4<= level3 & (7 downto 0 => '0') when ps(3)= '1' else     (7 downto 0 => '0') & level3;
   level5<= level4 & (15 downto 0 => '0') when ps(4)= '1' else     (15 downto 0 => '0') & level4;
   level6<= level5 & (31 downto 0 => '0') when ps(5)= '1' else     (31 downto 0 => '0') & level5;
   level7<= level6 & (63 downto 0 => '0') when ps(6)= '1' else     (63 downto 0 => '0') & level6;
   R <= level7(127 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                        PositDecoder_65_7_comb_uid16
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Raul Murillo, 2019
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity PositDecoder_65_7_comb_uid16 is
   port ( Input : in  std_logic_vector(64 downto 0);
          Sign : out  std_logic;
          Reg : out  std_logic_vector(7 downto 0);
          Exp : out  std_logic_vector(6 downto 0);
          Frac : out  std_logic_vector(55 downto 0);
          z : out  std_logic;
          inf : out  std_logic   );
end entity;

architecture arch of PositDecoder_65_7_comb_uid16 is
   component LZOC_64_comb_uid18 is
      port ( I : in  std_logic_vector(63 downto 0);
             OZB : in  std_logic;
             O : out  std_logic_vector(6 downto 0)   );
   end component;

   component LeftShifter_64_by_max_64_comb_uid22 is
      port ( X : in  std_logic_vector(63 downto 0);
             S : in  std_logic_vector(6 downto 0);
             R : out  std_logic_vector(127 downto 0)   );
   end component;

signal nzero :  std_logic;
signal my_sign :  std_logic;
signal rep_sign :  std_logic_vector(63 downto 0);
signal twos :  std_logic_vector(63 downto 0);
signal rc :  std_logic;
signal rep_rc :  std_logic_vector(63 downto 0);
signal inv :  std_logic_vector(63 downto 0);
signal zero_var :  std_logic;
signal zc :  std_logic_vector(6 downto 0);
signal zc_sub :  std_logic_vector(6 downto 0);
signal shifted_twos :  std_logic_vector(127 downto 0);
signal tmp :  std_logic_vector(61 downto 0);
begin
-------------------------------- Special Cases --------------------------------
   nzero <= '0' when Input(63 downto 0) = 0 else '1';
   -- 1 if Input is zero
   z <= Input(64) NOR nzero;
   -- 1 if Input is infinity
   inf <= Input(64) AND (NOT nzero);
------------------------------- Extract Sign bit -------------------------------
   my_sign <= Input(64);
   Sign <= my_sign;
--------------------------- 2's Complement of Input ---------------------------
   rep_sign <= (others => my_sign);
   twos <= (rep_sign XOR Input(63 downto 0)) + my_sign;
   rc <= twos(63);
------------------------ Count leading zeros of regime ------------------------
   rep_rc <= (others => rc);
   -- Invert 2's
   inv <= rep_rc XOR twos;
   zero_var <= '0';
   LZOC_Component: LZOC_64_comb_uid18
      port map ( I => inv,
                 O => zc,
                 OZB => zero_var);
----------------------------- Shift out the regime -----------------------------
   zc_sub <= zc - 1;
   LeftShifterComponent: LeftShifter_64_by_max_64_comb_uid22
      port map ( R => shifted_twos,
                 S => zc_sub,
                 X => twos);
   tmp <= shifted_twos(61 downto 0);
------------------------ Extract fraction and exponent ------------------------
   Frac <= nzero & tmp(54 downto 0);
   Exp <= tmp(61 downto 55);
-------------------------------- Select regime --------------------------------
   Reg <= '0' & zc_sub when rc = '1' else NOT('0' & zc) + 1;
end architecture;

--------------------------------------------------------------------------------
--                          IntAdder_113_f400_uid580
--                   (IntAdderAlternative_113_comb_uid584)
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2010)
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity IntAdder_113_f400_uid580 is
   port ( X : in  std_logic_vector(112 downto 0);
          Y : in  std_logic_vector(112 downto 0);
          Cin : in  std_logic;
          R : out  std_logic_vector(112 downto 0)   );
end entity;

architecture arch of IntAdder_113_f400_uid580 is
begin
   --Alternative
    R <= X + Y + Cin;
end architecture;

--------------------------------------------------------------------------------
--            IntMultiplier_UsingDSP_56_56_112_unsigned_comb_uid28
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Florent de Dinechin, Kinga Illyes, Bogdan Popa, Bogdan Pasca, 2012
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library std;
use std.textio.all;
library work;

entity IntMultiplier_UsingDSP_56_56_112_unsigned_comb_uid28 is
   port ( X : in  std_logic_vector(55 downto 0);
          Y : in  std_logic_vector(55 downto 0);
          R : out  std_logic_vector(111 downto 0)   );
end entity;

architecture arch of IntMultiplier_UsingDSP_56_56_112_unsigned_comb_uid28 is
   component IntAdder_113_f400_uid580 is
      port ( X : in  std_logic_vector(112 downto 0);
             Y : in  std_logic_vector(112 downto 0);
             Cin : in  std_logic;
             R : out  std_logic_vector(112 downto 0)   );
   end component;

   component SmallMultTableP3x3r6XuYu_comb_uid33 is
      port ( X : in  std_logic_vector(5 downto 0);
             Y : out  std_logic_vector(5 downto 0)   );
   end component;

   component SmallMultTableP3x3r6XuYu_comb_uid68 is
      port ( X : in  std_logic_vector(5 downto 0);
             Y : out  std_logic_vector(5 downto 0)   );
   end component;

   component SmallMultTableP3x3r6XuYu_comb_uid103 is
      port ( X : in  std_logic_vector(5 downto 0);
             Y : out  std_logic_vector(5 downto 0)   );
   end component;

   component Compressor_6_3 is
      port ( X0 : in  std_logic_vector(5 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_14_3 is
      port ( X0 : in  std_logic_vector(3 downto 0);
             X1 : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_5_3 is
      port ( X0 : in  std_logic_vector(4 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_4_3 is
      port ( X0 : in  std_logic_vector(3 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_23_3 is
      port ( X0 : in  std_logic_vector(2 downto 0);
             X1 : in  std_logic_vector(1 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_13_3 is
      port ( X0 : in  std_logic_vector(2 downto 0);
             X1 : in  std_logic_vector(0 downto 0);
             R : out  std_logic_vector(2 downto 0)   );
   end component;

   component Compressor_3_2 is
      port ( X0 : in  std_logic_vector(2 downto 0);
             R : out  std_logic_vector(1 downto 0)   );
   end component;

signal XX_m29 :  std_logic_vector(55 downto 0);
signal YY_m29 :  std_logic_vector(55 downto 0);
signal Xp_m29b31 :  std_logic_vector(23 downto 0);
signal Yp_m29b31 :  std_logic_vector(5 downto 0);
signal x_m29b31_0 :  std_logic_vector(2 downto 0);
signal x_m29b31_1 :  std_logic_vector(2 downto 0);
signal x_m29b31_2 :  std_logic_vector(2 downto 0);
signal x_m29b31_3 :  std_logic_vector(2 downto 0);
signal x_m29b31_4 :  std_logic_vector(2 downto 0);
signal x_m29b31_5 :  std_logic_vector(2 downto 0);
signal x_m29b31_6 :  std_logic_vector(2 downto 0);
signal x_m29b31_7 :  std_logic_vector(2 downto 0);
signal y_m29b31_0 :  std_logic_vector(2 downto 0);
signal y_m29b31_1 :  std_logic_vector(2 downto 0);
signal Y0X0_31_m29 :  std_logic_vector(5 downto 0);
signal PP31X0Y0_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w32_0 :  std_logic;
signal heap_bh30_w33_0 :  std_logic;
signal heap_bh30_w34_0 :  std_logic;
signal heap_bh30_w35_0 :  std_logic;
signal heap_bh30_w36_0 :  std_logic;
signal Y0X1_31_m29 :  std_logic_vector(5 downto 0);
signal PP31X1Y0_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w35_1 :  std_logic;
signal heap_bh30_w36_1 :  std_logic;
signal heap_bh30_w37_0 :  std_logic;
signal heap_bh30_w38_0 :  std_logic;
signal heap_bh30_w39_0 :  std_logic;
signal Y0X2_31_m29 :  std_logic_vector(5 downto 0);
signal PP31X2Y0_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w38_1 :  std_logic;
signal heap_bh30_w39_1 :  std_logic;
signal heap_bh30_w40_0 :  std_logic;
signal heap_bh30_w41_0 :  std_logic;
signal heap_bh30_w42_0 :  std_logic;
signal Y0X3_31_m29 :  std_logic_vector(5 downto 0);
signal PP31X3Y0_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w41_1 :  std_logic;
signal heap_bh30_w42_1 :  std_logic;
signal heap_bh30_w43_0 :  std_logic;
signal heap_bh30_w44_0 :  std_logic;
signal heap_bh30_w45_0 :  std_logic;
signal Y0X4_31_m29 :  std_logic_vector(5 downto 0);
signal PP31X4Y0_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w44_1 :  std_logic;
signal heap_bh30_w45_1 :  std_logic;
signal heap_bh30_w46_0 :  std_logic;
signal heap_bh30_w47_0 :  std_logic;
signal heap_bh30_w48_0 :  std_logic;
signal Y0X5_31_m29 :  std_logic_vector(5 downto 0);
signal PP31X5Y0_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w47_1 :  std_logic;
signal heap_bh30_w48_1 :  std_logic;
signal heap_bh30_w49_0 :  std_logic;
signal heap_bh30_w50_0 :  std_logic;
signal heap_bh30_w51_0 :  std_logic;
signal Y0X6_31_m29 :  std_logic_vector(5 downto 0);
signal PP31X6Y0_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w50_1 :  std_logic;
signal heap_bh30_w51_1 :  std_logic;
signal heap_bh30_w52_0 :  std_logic;
signal heap_bh30_w53_0 :  std_logic;
signal heap_bh30_w54_0 :  std_logic;
signal Y0X7_31_m29 :  std_logic_vector(5 downto 0);
signal PP31X7Y0_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w53_1 :  std_logic;
signal heap_bh30_w54_1 :  std_logic;
signal heap_bh30_w55_0 :  std_logic;
signal heap_bh30_w56_0 :  std_logic;
signal heap_bh30_w57_0 :  std_logic;
signal Y1X0_31_m29 :  std_logic_vector(5 downto 0);
signal PP31X0Y1_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w34_1 :  std_logic;
signal heap_bh30_w35_2 :  std_logic;
signal heap_bh30_w36_2 :  std_logic;
signal heap_bh30_w37_1 :  std_logic;
signal heap_bh30_w38_2 :  std_logic;
signal heap_bh30_w39_2 :  std_logic;
signal Y1X1_31_m29 :  std_logic_vector(5 downto 0);
signal PP31X1Y1_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w37_2 :  std_logic;
signal heap_bh30_w38_3 :  std_logic;
signal heap_bh30_w39_3 :  std_logic;
signal heap_bh30_w40_1 :  std_logic;
signal heap_bh30_w41_2 :  std_logic;
signal heap_bh30_w42_2 :  std_logic;
signal Y1X2_31_m29 :  std_logic_vector(5 downto 0);
signal PP31X2Y1_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w40_2 :  std_logic;
signal heap_bh30_w41_3 :  std_logic;
signal heap_bh30_w42_3 :  std_logic;
signal heap_bh30_w43_1 :  std_logic;
signal heap_bh30_w44_2 :  std_logic;
signal heap_bh30_w45_2 :  std_logic;
signal Y1X3_31_m29 :  std_logic_vector(5 downto 0);
signal PP31X3Y1_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w43_2 :  std_logic;
signal heap_bh30_w44_3 :  std_logic;
signal heap_bh30_w45_3 :  std_logic;
signal heap_bh30_w46_1 :  std_logic;
signal heap_bh30_w47_2 :  std_logic;
signal heap_bh30_w48_2 :  std_logic;
signal Y1X4_31_m29 :  std_logic_vector(5 downto 0);
signal PP31X4Y1_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w46_2 :  std_logic;
signal heap_bh30_w47_3 :  std_logic;
signal heap_bh30_w48_3 :  std_logic;
signal heap_bh30_w49_1 :  std_logic;
signal heap_bh30_w50_2 :  std_logic;
signal heap_bh30_w51_2 :  std_logic;
signal Y1X5_31_m29 :  std_logic_vector(5 downto 0);
signal PP31X5Y1_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w49_2 :  std_logic;
signal heap_bh30_w50_3 :  std_logic;
signal heap_bh30_w51_3 :  std_logic;
signal heap_bh30_w52_1 :  std_logic;
signal heap_bh30_w53_2 :  std_logic;
signal heap_bh30_w54_2 :  std_logic;
signal Y1X6_31_m29 :  std_logic_vector(5 downto 0);
signal PP31X6Y1_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w52_2 :  std_logic;
signal heap_bh30_w53_3 :  std_logic;
signal heap_bh30_w54_3 :  std_logic;
signal heap_bh30_w55_1 :  std_logic;
signal heap_bh30_w56_1 :  std_logic;
signal heap_bh30_w57_1 :  std_logic;
signal Y1X7_31_m29 :  std_logic_vector(5 downto 0);
signal PP31X7Y1_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w55_2 :  std_logic;
signal heap_bh30_w56_2 :  std_logic;
signal heap_bh30_w57_2 :  std_logic;
signal heap_bh30_w58_0 :  std_logic;
signal heap_bh30_w59_0 :  std_logic;
signal heap_bh30_w60_0 :  std_logic;
signal Xp_m29b66 :  std_logic_vector(23 downto 0);
signal Yp_m29b66 :  std_logic_vector(5 downto 0);
signal x_m29b66_0 :  std_logic_vector(2 downto 0);
signal x_m29b66_1 :  std_logic_vector(2 downto 0);
signal x_m29b66_2 :  std_logic_vector(2 downto 0);
signal x_m29b66_3 :  std_logic_vector(2 downto 0);
signal x_m29b66_4 :  std_logic_vector(2 downto 0);
signal x_m29b66_5 :  std_logic_vector(2 downto 0);
signal x_m29b66_6 :  std_logic_vector(2 downto 0);
signal x_m29b66_7 :  std_logic_vector(2 downto 0);
signal y_m29b66_0 :  std_logic_vector(2 downto 0);
signal y_m29b66_1 :  std_logic_vector(2 downto 0);
signal Y0X0_66_m29 :  std_logic_vector(5 downto 0);
signal PP66X0Y0_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w8_0 :  std_logic;
signal heap_bh30_w9_0 :  std_logic;
signal heap_bh30_w10_0 :  std_logic;
signal heap_bh30_w11_0 :  std_logic;
signal heap_bh30_w12_0 :  std_logic;
signal Y0X1_66_m29 :  std_logic_vector(5 downto 0);
signal PP66X1Y0_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w11_1 :  std_logic;
signal heap_bh30_w12_1 :  std_logic;
signal heap_bh30_w13_0 :  std_logic;
signal heap_bh30_w14_0 :  std_logic;
signal heap_bh30_w15_0 :  std_logic;
signal Y0X2_66_m29 :  std_logic_vector(5 downto 0);
signal PP66X2Y0_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w14_1 :  std_logic;
signal heap_bh30_w15_1 :  std_logic;
signal heap_bh30_w16_0 :  std_logic;
signal heap_bh30_w17_0 :  std_logic;
signal heap_bh30_w18_0 :  std_logic;
signal Y0X3_66_m29 :  std_logic_vector(5 downto 0);
signal PP66X3Y0_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w17_1 :  std_logic;
signal heap_bh30_w18_1 :  std_logic;
signal heap_bh30_w19_0 :  std_logic;
signal heap_bh30_w20_0 :  std_logic;
signal heap_bh30_w21_0 :  std_logic;
signal Y0X4_66_m29 :  std_logic_vector(5 downto 0);
signal PP66X4Y0_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w20_1 :  std_logic;
signal heap_bh30_w21_1 :  std_logic;
signal heap_bh30_w22_0 :  std_logic;
signal heap_bh30_w23_0 :  std_logic;
signal heap_bh30_w24_0 :  std_logic;
signal Y0X5_66_m29 :  std_logic_vector(5 downto 0);
signal PP66X5Y0_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w23_1 :  std_logic;
signal heap_bh30_w24_1 :  std_logic;
signal heap_bh30_w25_0 :  std_logic;
signal heap_bh30_w26_0 :  std_logic;
signal heap_bh30_w27_0 :  std_logic;
signal Y0X6_66_m29 :  std_logic_vector(5 downto 0);
signal PP66X6Y0_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w26_1 :  std_logic;
signal heap_bh30_w27_1 :  std_logic;
signal heap_bh30_w28_0 :  std_logic;
signal heap_bh30_w29_0 :  std_logic;
signal heap_bh30_w30_0 :  std_logic;
signal Y0X7_66_m29 :  std_logic_vector(5 downto 0);
signal PP66X7Y0_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w29_1 :  std_logic;
signal heap_bh30_w30_1 :  std_logic;
signal heap_bh30_w31_0 :  std_logic;
signal heap_bh30_w32_1 :  std_logic;
signal heap_bh30_w33_1 :  std_logic;
signal Y1X0_66_m29 :  std_logic_vector(5 downto 0);
signal PP66X0Y1_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w10_1 :  std_logic;
signal heap_bh30_w11_2 :  std_logic;
signal heap_bh30_w12_2 :  std_logic;
signal heap_bh30_w13_1 :  std_logic;
signal heap_bh30_w14_2 :  std_logic;
signal heap_bh30_w15_2 :  std_logic;
signal Y1X1_66_m29 :  std_logic_vector(5 downto 0);
signal PP66X1Y1_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w13_2 :  std_logic;
signal heap_bh30_w14_3 :  std_logic;
signal heap_bh30_w15_3 :  std_logic;
signal heap_bh30_w16_1 :  std_logic;
signal heap_bh30_w17_2 :  std_logic;
signal heap_bh30_w18_2 :  std_logic;
signal Y1X2_66_m29 :  std_logic_vector(5 downto 0);
signal PP66X2Y1_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w16_2 :  std_logic;
signal heap_bh30_w17_3 :  std_logic;
signal heap_bh30_w18_3 :  std_logic;
signal heap_bh30_w19_1 :  std_logic;
signal heap_bh30_w20_2 :  std_logic;
signal heap_bh30_w21_2 :  std_logic;
signal Y1X3_66_m29 :  std_logic_vector(5 downto 0);
signal PP66X3Y1_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w19_2 :  std_logic;
signal heap_bh30_w20_3 :  std_logic;
signal heap_bh30_w21_3 :  std_logic;
signal heap_bh30_w22_1 :  std_logic;
signal heap_bh30_w23_2 :  std_logic;
signal heap_bh30_w24_2 :  std_logic;
signal Y1X4_66_m29 :  std_logic_vector(5 downto 0);
signal PP66X4Y1_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w22_2 :  std_logic;
signal heap_bh30_w23_3 :  std_logic;
signal heap_bh30_w24_3 :  std_logic;
signal heap_bh30_w25_1 :  std_logic;
signal heap_bh30_w26_2 :  std_logic;
signal heap_bh30_w27_2 :  std_logic;
signal Y1X5_66_m29 :  std_logic_vector(5 downto 0);
signal PP66X5Y1_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w25_2 :  std_logic;
signal heap_bh30_w26_3 :  std_logic;
signal heap_bh30_w27_3 :  std_logic;
signal heap_bh30_w28_1 :  std_logic;
signal heap_bh30_w29_2 :  std_logic;
signal heap_bh30_w30_2 :  std_logic;
signal Y1X6_66_m29 :  std_logic_vector(5 downto 0);
signal PP66X6Y1_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w28_2 :  std_logic;
signal heap_bh30_w29_3 :  std_logic;
signal heap_bh30_w30_3 :  std_logic;
signal heap_bh30_w31_1 :  std_logic;
signal heap_bh30_w32_2 :  std_logic;
signal heap_bh30_w33_2 :  std_logic;
signal Y1X7_66_m29 :  std_logic_vector(5 downto 0);
signal PP66X7Y1_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w31_2 :  std_logic;
signal heap_bh30_w32_3 :  std_logic;
signal heap_bh30_w33_3 :  std_logic;
signal heap_bh30_w34_2 :  std_logic;
signal heap_bh30_w35_3 :  std_logic;
signal heap_bh30_w36_3 :  std_logic;
signal Xp_m29b101 :  std_logic_vector(8 downto 0);
signal Yp_m29b101 :  std_logic_vector(5 downto 0);
signal x_m29b101_0 :  std_logic_vector(2 downto 0);
signal x_m29b101_1 :  std_logic_vector(2 downto 0);
signal x_m29b101_2 :  std_logic_vector(2 downto 0);
signal y_m29b101_0 :  std_logic_vector(2 downto 0);
signal y_m29b101_1 :  std_logic_vector(2 downto 0);
signal Y0X0_101_m29 :  std_logic_vector(5 downto 0);
signal PP101X0Y0_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w0_0 :  std_logic;
signal heap_bh30_w1_0 :  std_logic;
signal heap_bh30_w2_0 :  std_logic;
signal heap_bh30_w3_0 :  std_logic;
signal Y0X1_101_m29 :  std_logic_vector(5 downto 0);
signal PP101X1Y0_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w2_1 :  std_logic;
signal heap_bh30_w3_1 :  std_logic;
signal heap_bh30_w4_0 :  std_logic;
signal heap_bh30_w5_0 :  std_logic;
signal heap_bh30_w6_0 :  std_logic;
signal Y0X2_101_m29 :  std_logic_vector(5 downto 0);
signal PP101X2Y0_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w5_1 :  std_logic;
signal heap_bh30_w6_1 :  std_logic;
signal heap_bh30_w7_0 :  std_logic;
signal heap_bh30_w8_1 :  std_logic;
signal heap_bh30_w9_1 :  std_logic;
signal Y1X0_101_m29 :  std_logic_vector(5 downto 0);
signal PP101X0Y1_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w2_2 :  std_logic;
signal heap_bh30_w3_2 :  std_logic;
signal heap_bh30_w4_1 :  std_logic;
signal heap_bh30_w5_2 :  std_logic;
signal heap_bh30_w6_2 :  std_logic;
signal Y1X1_101_m29 :  std_logic_vector(5 downto 0);
signal PP101X1Y1_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w4_2 :  std_logic;
signal heap_bh30_w5_3 :  std_logic;
signal heap_bh30_w6_3 :  std_logic;
signal heap_bh30_w7_1 :  std_logic;
signal heap_bh30_w8_2 :  std_logic;
signal heap_bh30_w9_2 :  std_logic;
signal Y1X2_101_m29 :  std_logic_vector(5 downto 0);
signal PP101X2Y1_m29 :  std_logic_vector(5 downto 0);
signal heap_bh30_w7_2 :  std_logic;
signal heap_bh30_w8_3 :  std_logic;
signal heap_bh30_w9_3 :  std_logic;
signal heap_bh30_w10_2 :  std_logic;
signal heap_bh30_w11_3 :  std_logic;
signal heap_bh30_w12_3 :  std_logic;
signal DSP_bh30_ch0_0 :  std_logic_vector(40 downto 0);
signal heap_bh30_w111_0 :  std_logic;
signal heap_bh30_w110_0 :  std_logic;
signal heap_bh30_w109_0 :  std_logic;
signal heap_bh30_w108_0 :  std_logic;
signal heap_bh30_w107_0 :  std_logic;
signal heap_bh30_w106_0 :  std_logic;
signal heap_bh30_w105_0 :  std_logic;
signal heap_bh30_w104_0 :  std_logic;
signal heap_bh30_w103_0 :  std_logic;
signal heap_bh30_w102_0 :  std_logic;
signal heap_bh30_w101_0 :  std_logic;
signal heap_bh30_w100_0 :  std_logic;
signal heap_bh30_w99_0 :  std_logic;
signal heap_bh30_w98_0 :  std_logic;
signal heap_bh30_w97_0 :  std_logic;
signal heap_bh30_w96_0 :  std_logic;
signal heap_bh30_w95_0 :  std_logic;
signal heap_bh30_w94_0 :  std_logic;
signal heap_bh30_w93_0 :  std_logic;
signal heap_bh30_w92_0 :  std_logic;
signal heap_bh30_w91_0 :  std_logic;
signal heap_bh30_w90_0 :  std_logic;
signal heap_bh30_w89_0 :  std_logic;
signal heap_bh30_w88_0 :  std_logic;
signal heap_bh30_w87_0 :  std_logic;
signal heap_bh30_w86_0 :  std_logic;
signal heap_bh30_w85_0 :  std_logic;
signal heap_bh30_w84_0 :  std_logic;
signal heap_bh30_w83_0 :  std_logic;
signal heap_bh30_w82_0 :  std_logic;
signal heap_bh30_w81_0 :  std_logic;
signal heap_bh30_w80_0 :  std_logic;
signal heap_bh30_w79_0 :  std_logic;
signal heap_bh30_w78_0 :  std_logic;
signal heap_bh30_w77_0 :  std_logic;
signal heap_bh30_w76_0 :  std_logic;
signal heap_bh30_w75_0 :  std_logic;
signal heap_bh30_w74_0 :  std_logic;
signal heap_bh30_w73_0 :  std_logic;
signal heap_bh30_w72_0 :  std_logic;
signal heap_bh30_w71_0 :  std_logic;
signal DSP_bh30_ch1_0 :  std_logic_vector(40 downto 0);
signal heap_bh30_w87_1 :  std_logic;
signal heap_bh30_w86_1 :  std_logic;
signal heap_bh30_w85_1 :  std_logic;
signal heap_bh30_w84_1 :  std_logic;
signal heap_bh30_w83_1 :  std_logic;
signal heap_bh30_w82_1 :  std_logic;
signal heap_bh30_w81_1 :  std_logic;
signal heap_bh30_w80_1 :  std_logic;
signal heap_bh30_w79_1 :  std_logic;
signal heap_bh30_w78_1 :  std_logic;
signal heap_bh30_w77_1 :  std_logic;
signal heap_bh30_w76_1 :  std_logic;
signal heap_bh30_w75_1 :  std_logic;
signal heap_bh30_w74_1 :  std_logic;
signal heap_bh30_w73_1 :  std_logic;
signal heap_bh30_w72_1 :  std_logic;
signal heap_bh30_w71_1 :  std_logic;
signal heap_bh30_w70_0 :  std_logic;
signal heap_bh30_w69_0 :  std_logic;
signal heap_bh30_w68_0 :  std_logic;
signal heap_bh30_w67_0 :  std_logic;
signal heap_bh30_w66_0 :  std_logic;
signal heap_bh30_w65_0 :  std_logic;
signal heap_bh30_w64_0 :  std_logic;
signal heap_bh30_w63_0 :  std_logic;
signal heap_bh30_w62_0 :  std_logic;
signal heap_bh30_w61_0 :  std_logic;
signal heap_bh30_w60_1 :  std_logic;
signal heap_bh30_w59_1 :  std_logic;
signal heap_bh30_w58_1 :  std_logic;
signal heap_bh30_w57_3 :  std_logic;
signal heap_bh30_w56_3 :  std_logic;
signal heap_bh30_w55_3 :  std_logic;
signal heap_bh30_w54_4 :  std_logic;
signal heap_bh30_w53_4 :  std_logic;
signal heap_bh30_w52_3 :  std_logic;
signal heap_bh30_w51_4 :  std_logic;
signal heap_bh30_w50_4 :  std_logic;
signal heap_bh30_w49_3 :  std_logic;
signal heap_bh30_w48_4 :  std_logic;
signal heap_bh30_w47_4 :  std_logic;
signal DSP_bh30_ch2_0 :  std_logic_vector(40 downto 0);
signal heap_bh30_w63_1 :  std_logic;
signal heap_bh30_w62_1 :  std_logic;
signal heap_bh30_w61_1 :  std_logic;
signal heap_bh30_w60_2 :  std_logic;
signal heap_bh30_w59_2 :  std_logic;
signal heap_bh30_w58_2 :  std_logic;
signal heap_bh30_w57_4 :  std_logic;
signal heap_bh30_w56_4 :  std_logic;
signal heap_bh30_w55_4 :  std_logic;
signal heap_bh30_w54_5 :  std_logic;
signal heap_bh30_w53_5 :  std_logic;
signal heap_bh30_w52_4 :  std_logic;
signal heap_bh30_w51_5 :  std_logic;
signal heap_bh30_w50_5 :  std_logic;
signal heap_bh30_w49_4 :  std_logic;
signal heap_bh30_w48_5 :  std_logic;
signal heap_bh30_w47_5 :  std_logic;
signal heap_bh30_w46_3 :  std_logic;
signal heap_bh30_w45_4 :  std_logic;
signal heap_bh30_w44_4 :  std_logic;
signal heap_bh30_w43_3 :  std_logic;
signal heap_bh30_w42_4 :  std_logic;
signal heap_bh30_w41_4 :  std_logic;
signal heap_bh30_w40_3 :  std_logic;
signal heap_bh30_w39_4 :  std_logic;
signal heap_bh30_w38_4 :  std_logic;
signal heap_bh30_w37_3 :  std_logic;
signal heap_bh30_w36_4 :  std_logic;
signal heap_bh30_w35_4 :  std_logic;
signal heap_bh30_w34_3 :  std_logic;
signal heap_bh30_w33_4 :  std_logic;
signal heap_bh30_w32_4 :  std_logic;
signal heap_bh30_w31_3 :  std_logic;
signal heap_bh30_w30_4 :  std_logic;
signal heap_bh30_w29_4 :  std_logic;
signal heap_bh30_w28_3 :  std_logic;
signal heap_bh30_w27_4 :  std_logic;
signal heap_bh30_w26_4 :  std_logic;
signal heap_bh30_w25_3 :  std_logic;
signal heap_bh30_w24_4 :  std_logic;
signal heap_bh30_w23_4 :  std_logic;
signal DSP_bh30_ch3_0 :  std_logic_vector(40 downto 0);
signal heap_bh30_w94_1 :  std_logic;
signal heap_bh30_w93_1 :  std_logic;
signal heap_bh30_w92_1 :  std_logic;
signal heap_bh30_w91_1 :  std_logic;
signal heap_bh30_w90_1 :  std_logic;
signal heap_bh30_w89_1 :  std_logic;
signal heap_bh30_w88_1 :  std_logic;
signal heap_bh30_w87_2 :  std_logic;
signal heap_bh30_w86_2 :  std_logic;
signal heap_bh30_w85_2 :  std_logic;
signal heap_bh30_w84_2 :  std_logic;
signal heap_bh30_w83_2 :  std_logic;
signal heap_bh30_w82_2 :  std_logic;
signal heap_bh30_w81_2 :  std_logic;
signal heap_bh30_w80_2 :  std_logic;
signal heap_bh30_w79_2 :  std_logic;
signal heap_bh30_w78_2 :  std_logic;
signal heap_bh30_w77_2 :  std_logic;
signal heap_bh30_w76_2 :  std_logic;
signal heap_bh30_w75_2 :  std_logic;
signal heap_bh30_w74_2 :  std_logic;
signal heap_bh30_w73_2 :  std_logic;
signal heap_bh30_w72_2 :  std_logic;
signal heap_bh30_w71_2 :  std_logic;
signal heap_bh30_w70_1 :  std_logic;
signal heap_bh30_w69_1 :  std_logic;
signal heap_bh30_w68_1 :  std_logic;
signal heap_bh30_w67_1 :  std_logic;
signal heap_bh30_w66_1 :  std_logic;
signal heap_bh30_w65_1 :  std_logic;
signal heap_bh30_w64_1 :  std_logic;
signal heap_bh30_w63_2 :  std_logic;
signal heap_bh30_w62_2 :  std_logic;
signal heap_bh30_w61_2 :  std_logic;
signal heap_bh30_w60_3 :  std_logic;
signal heap_bh30_w59_3 :  std_logic;
signal heap_bh30_w58_3 :  std_logic;
signal heap_bh30_w57_5 :  std_logic;
signal heap_bh30_w56_5 :  std_logic;
signal heap_bh30_w55_5 :  std_logic;
signal heap_bh30_w54_6 :  std_logic;
signal DSP_bh30_ch4_0 :  std_logic_vector(40 downto 0);
signal heap_bh30_w70_2 :  std_logic;
signal heap_bh30_w69_2 :  std_logic;
signal heap_bh30_w68_2 :  std_logic;
signal heap_bh30_w67_2 :  std_logic;
signal heap_bh30_w66_2 :  std_logic;
signal heap_bh30_w65_2 :  std_logic;
signal heap_bh30_w64_2 :  std_logic;
signal heap_bh30_w63_3 :  std_logic;
signal heap_bh30_w62_3 :  std_logic;
signal heap_bh30_w61_3 :  std_logic;
signal heap_bh30_w60_4 :  std_logic;
signal heap_bh30_w59_4 :  std_logic;
signal heap_bh30_w58_4 :  std_logic;
signal heap_bh30_w57_6 :  std_logic;
signal heap_bh30_w56_6 :  std_logic;
signal heap_bh30_w55_6 :  std_logic;
signal heap_bh30_w54_7 :  std_logic;
signal heap_bh30_w53_6 :  std_logic;
signal heap_bh30_w52_5 :  std_logic;
signal heap_bh30_w51_6 :  std_logic;
signal heap_bh30_w50_6 :  std_logic;
signal heap_bh30_w49_5 :  std_logic;
signal heap_bh30_w48_6 :  std_logic;
signal heap_bh30_w47_6 :  std_logic;
signal heap_bh30_w46_4 :  std_logic;
signal heap_bh30_w45_5 :  std_logic;
signal heap_bh30_w44_5 :  std_logic;
signal heap_bh30_w43_4 :  std_logic;
signal heap_bh30_w42_5 :  std_logic;
signal heap_bh30_w41_5 :  std_logic;
signal heap_bh30_w40_4 :  std_logic;
signal heap_bh30_w39_5 :  std_logic;
signal heap_bh30_w38_5 :  std_logic;
signal heap_bh30_w37_4 :  std_logic;
signal heap_bh30_w36_5 :  std_logic;
signal heap_bh30_w35_5 :  std_logic;
signal heap_bh30_w34_4 :  std_logic;
signal heap_bh30_w33_5 :  std_logic;
signal heap_bh30_w32_5 :  std_logic;
signal heap_bh30_w31_4 :  std_logic;
signal heap_bh30_w30_5 :  std_logic;
signal DSP_bh30_ch5_0 :  std_logic_vector(40 downto 0);
signal heap_bh30_w46_5 :  std_logic;
signal heap_bh30_w45_6 :  std_logic;
signal heap_bh30_w44_6 :  std_logic;
signal heap_bh30_w43_5 :  std_logic;
signal heap_bh30_w42_6 :  std_logic;
signal heap_bh30_w41_6 :  std_logic;
signal heap_bh30_w40_5 :  std_logic;
signal heap_bh30_w39_6 :  std_logic;
signal heap_bh30_w38_6 :  std_logic;
signal heap_bh30_w37_5 :  std_logic;
signal heap_bh30_w36_6 :  std_logic;
signal heap_bh30_w35_6 :  std_logic;
signal heap_bh30_w34_5 :  std_logic;
signal heap_bh30_w33_6 :  std_logic;
signal heap_bh30_w32_6 :  std_logic;
signal heap_bh30_w31_5 :  std_logic;
signal heap_bh30_w30_6 :  std_logic;
signal heap_bh30_w29_5 :  std_logic;
signal heap_bh30_w28_4 :  std_logic;
signal heap_bh30_w27_5 :  std_logic;
signal heap_bh30_w26_5 :  std_logic;
signal heap_bh30_w25_4 :  std_logic;
signal heap_bh30_w24_5 :  std_logic;
signal heap_bh30_w23_5 :  std_logic;
signal heap_bh30_w22_3 :  std_logic;
signal heap_bh30_w21_4 :  std_logic;
signal heap_bh30_w20_4 :  std_logic;
signal heap_bh30_w19_3 :  std_logic;
signal heap_bh30_w18_4 :  std_logic;
signal heap_bh30_w17_4 :  std_logic;
signal heap_bh30_w16_3 :  std_logic;
signal heap_bh30_w15_4 :  std_logic;
signal heap_bh30_w14_4 :  std_logic;
signal heap_bh30_w13_3 :  std_logic;
signal heap_bh30_w12_4 :  std_logic;
signal heap_bh30_w11_4 :  std_logic;
signal heap_bh30_w10_3 :  std_logic;
signal heap_bh30_w9_4 :  std_logic;
signal heap_bh30_w8_4 :  std_logic;
signal heap_bh30_w7_3 :  std_logic;
signal heap_bh30_w6_4 :  std_logic;
signal DSP_bh30_ch6_0 :  std_logic_vector(40 downto 0);
signal heap_bh30_w77_3 :  std_logic;
signal heap_bh30_w76_3 :  std_logic;
signal heap_bh30_w75_3 :  std_logic;
signal heap_bh30_w74_3 :  std_logic;
signal heap_bh30_w73_3 :  std_logic;
signal heap_bh30_w72_3 :  std_logic;
signal heap_bh30_w71_3 :  std_logic;
signal heap_bh30_w70_3 :  std_logic;
signal heap_bh30_w69_3 :  std_logic;
signal heap_bh30_w68_3 :  std_logic;
signal heap_bh30_w67_3 :  std_logic;
signal heap_bh30_w66_3 :  std_logic;
signal heap_bh30_w65_3 :  std_logic;
signal heap_bh30_w64_3 :  std_logic;
signal heap_bh30_w63_4 :  std_logic;
signal heap_bh30_w62_4 :  std_logic;
signal heap_bh30_w61_4 :  std_logic;
signal heap_bh30_w60_5 :  std_logic;
signal heap_bh30_w59_5 :  std_logic;
signal heap_bh30_w58_5 :  std_logic;
signal heap_bh30_w57_7 :  std_logic;
signal heap_bh30_w56_7 :  std_logic;
signal heap_bh30_w55_7 :  std_logic;
signal heap_bh30_w54_8 :  std_logic;
signal heap_bh30_w53_7 :  std_logic;
signal heap_bh30_w52_6 :  std_logic;
signal heap_bh30_w51_7 :  std_logic;
signal heap_bh30_w50_7 :  std_logic;
signal heap_bh30_w49_6 :  std_logic;
signal heap_bh30_w48_7 :  std_logic;
signal heap_bh30_w47_7 :  std_logic;
signal heap_bh30_w46_6 :  std_logic;
signal heap_bh30_w45_7 :  std_logic;
signal heap_bh30_w44_7 :  std_logic;
signal heap_bh30_w43_6 :  std_logic;
signal heap_bh30_w42_7 :  std_logic;
signal heap_bh30_w41_7 :  std_logic;
signal heap_bh30_w40_6 :  std_logic;
signal heap_bh30_w39_7 :  std_logic;
signal heap_bh30_w38_7 :  std_logic;
signal heap_bh30_w37_6 :  std_logic;
signal DSP_bh30_ch7_0 :  std_logic_vector(40 downto 0);
signal heap_bh30_w53_8 :  std_logic;
signal heap_bh30_w52_7 :  std_logic;
signal heap_bh30_w51_8 :  std_logic;
signal heap_bh30_w50_8 :  std_logic;
signal heap_bh30_w49_7 :  std_logic;
signal heap_bh30_w48_8 :  std_logic;
signal heap_bh30_w47_8 :  std_logic;
signal heap_bh30_w46_7 :  std_logic;
signal heap_bh30_w45_8 :  std_logic;
signal heap_bh30_w44_8 :  std_logic;
signal heap_bh30_w43_7 :  std_logic;
signal heap_bh30_w42_8 :  std_logic;
signal heap_bh30_w41_8 :  std_logic;
signal heap_bh30_w40_7 :  std_logic;
signal heap_bh30_w39_8 :  std_logic;
signal heap_bh30_w38_8 :  std_logic;
signal heap_bh30_w37_7 :  std_logic;
signal heap_bh30_w36_7 :  std_logic;
signal heap_bh30_w35_7 :  std_logic;
signal heap_bh30_w34_6 :  std_logic;
signal heap_bh30_w33_7 :  std_logic;
signal heap_bh30_w32_7 :  std_logic;
signal heap_bh30_w31_6 :  std_logic;
signal heap_bh30_w30_7 :  std_logic;
signal heap_bh30_w29_6 :  std_logic;
signal heap_bh30_w28_5 :  std_logic;
signal heap_bh30_w27_6 :  std_logic;
signal heap_bh30_w26_6 :  std_logic;
signal heap_bh30_w25_5 :  std_logic;
signal heap_bh30_w24_6 :  std_logic;
signal heap_bh30_w23_6 :  std_logic;
signal heap_bh30_w22_4 :  std_logic;
signal heap_bh30_w21_5 :  std_logic;
signal heap_bh30_w20_5 :  std_logic;
signal heap_bh30_w19_4 :  std_logic;
signal heap_bh30_w18_5 :  std_logic;
signal heap_bh30_w17_5 :  std_logic;
signal heap_bh30_w16_4 :  std_logic;
signal heap_bh30_w15_5 :  std_logic;
signal heap_bh30_w14_5 :  std_logic;
signal heap_bh30_w13_4 :  std_logic;
signal DSP_bh30_ch8_0 :  std_logic_vector(40 downto 0);
signal heap_bh30_w29_7 :  std_logic;
signal heap_bh30_w28_6 :  std_logic;
signal heap_bh30_w27_7 :  std_logic;
signal heap_bh30_w26_7 :  std_logic;
signal heap_bh30_w25_6 :  std_logic;
signal heap_bh30_w24_7 :  std_logic;
signal heap_bh30_w23_7 :  std_logic;
signal heap_bh30_w22_5 :  std_logic;
signal heap_bh30_w21_6 :  std_logic;
signal heap_bh30_w20_6 :  std_logic;
signal heap_bh30_w19_5 :  std_logic;
signal heap_bh30_w18_6 :  std_logic;
signal heap_bh30_w17_6 :  std_logic;
signal heap_bh30_w16_5 :  std_logic;
signal heap_bh30_w15_6 :  std_logic;
signal heap_bh30_w14_6 :  std_logic;
signal heap_bh30_w13_5 :  std_logic;
signal heap_bh30_w12_5 :  std_logic;
signal heap_bh30_w11_5 :  std_logic;
signal heap_bh30_w10_4 :  std_logic;
signal heap_bh30_w9_5 :  std_logic;
signal heap_bh30_w8_5 :  std_logic;
signal heap_bh30_w7_4 :  std_logic;
signal heap_bh30_w6_5 :  std_logic;
signal heap_bh30_w5_4 :  std_logic;
signal heap_bh30_w4_3 :  std_logic;
signal heap_bh30_w3_3 :  std_logic;
signal heap_bh30_w2_3 :  std_logic;
signal heap_bh30_w1_1 :  std_logic;
signal heap_bh30_w0_1 :  std_logic;
signal CompressorIn_bh30_0_0 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_0_1 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_0_0 :  std_logic_vector(2 downto 0);
signal heap_bh30_w5_5 :  std_logic;
signal heap_bh30_w6_6 :  std_logic;
signal heap_bh30_w7_5 :  std_logic;
signal CompressorIn_bh30_1_2 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_1_3 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_1_1 :  std_logic_vector(2 downto 0);
signal heap_bh30_w8_6 :  std_logic;
signal heap_bh30_w9_6 :  std_logic;
signal heap_bh30_w10_5 :  std_logic;
signal CompressorIn_bh30_2_4 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_2_5 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_2_2 :  std_logic_vector(2 downto 0);
signal heap_bh30_w11_6 :  std_logic;
signal heap_bh30_w12_6 :  std_logic;
signal heap_bh30_w13_6 :  std_logic;
signal CompressorIn_bh30_3_6 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_3_7 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_3_3 :  std_logic_vector(2 downto 0);
signal heap_bh30_w14_7 :  std_logic;
signal heap_bh30_w15_7 :  std_logic;
signal heap_bh30_w16_6 :  std_logic;
signal CompressorIn_bh30_4_8 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_4_9 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_4_4 :  std_logic_vector(2 downto 0);
signal heap_bh30_w17_7 :  std_logic;
signal heap_bh30_w18_7 :  std_logic;
signal heap_bh30_w19_6 :  std_logic;
signal CompressorIn_bh30_5_10 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_5_11 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_5_5 :  std_logic_vector(2 downto 0);
signal heap_bh30_w20_7 :  std_logic;
signal heap_bh30_w21_7 :  std_logic;
signal heap_bh30_w22_6 :  std_logic;
signal CompressorIn_bh30_6_12 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_6_13 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_6_6 :  std_logic_vector(2 downto 0);
signal heap_bh30_w23_8 :  std_logic;
signal heap_bh30_w24_8 :  std_logic;
signal heap_bh30_w25_7 :  std_logic;
signal CompressorIn_bh30_7_14 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_7_15 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_7_7 :  std_logic_vector(2 downto 0);
signal heap_bh30_w26_8 :  std_logic;
signal heap_bh30_w27_8 :  std_logic;
signal heap_bh30_w28_7 :  std_logic;
signal CompressorIn_bh30_8_16 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_8_17 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_8_8 :  std_logic_vector(2 downto 0);
signal heap_bh30_w29_8 :  std_logic;
signal heap_bh30_w30_8 :  std_logic;
signal heap_bh30_w31_7 :  std_logic;
signal CompressorIn_bh30_9_18 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_9_19 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_9_9 :  std_logic_vector(2 downto 0);
signal heap_bh30_w32_8 :  std_logic;
signal heap_bh30_w33_8 :  std_logic;
signal heap_bh30_w34_7 :  std_logic;
signal CompressorIn_bh30_10_20 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_10_21 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_10_10 :  std_logic_vector(2 downto 0);
signal heap_bh30_w35_8 :  std_logic;
signal heap_bh30_w36_8 :  std_logic;
signal heap_bh30_w37_8 :  std_logic;
signal CompressorIn_bh30_11_22 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_11_23 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_11_11 :  std_logic_vector(2 downto 0);
signal heap_bh30_w38_9 :  std_logic;
signal heap_bh30_w39_9 :  std_logic;
signal heap_bh30_w40_8 :  std_logic;
signal CompressorIn_bh30_12_24 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_12_25 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_12_12 :  std_logic_vector(2 downto 0);
signal heap_bh30_w41_9 :  std_logic;
signal heap_bh30_w42_9 :  std_logic;
signal heap_bh30_w43_8 :  std_logic;
signal CompressorIn_bh30_13_26 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_13_27 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_13_13 :  std_logic_vector(2 downto 0);
signal heap_bh30_w44_9 :  std_logic;
signal heap_bh30_w45_9 :  std_logic;
signal heap_bh30_w46_8 :  std_logic;
signal CompressorIn_bh30_14_28 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_14_29 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_14_14 :  std_logic_vector(2 downto 0);
signal heap_bh30_w47_9 :  std_logic;
signal heap_bh30_w48_9 :  std_logic;
signal heap_bh30_w49_8 :  std_logic;
signal CompressorIn_bh30_15_30 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_15_31 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_15_15 :  std_logic_vector(2 downto 0);
signal heap_bh30_w50_9 :  std_logic;
signal heap_bh30_w51_9 :  std_logic;
signal heap_bh30_w52_8 :  std_logic;
signal CompressorIn_bh30_16_32 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_16_33 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_16_16 :  std_logic_vector(2 downto 0);
signal heap_bh30_w53_9 :  std_logic;
signal heap_bh30_w54_9 :  std_logic;
signal heap_bh30_w55_8 :  std_logic;
signal CompressorIn_bh30_17_34 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_17_35 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_17_17 :  std_logic_vector(2 downto 0);
signal heap_bh30_w2_4 :  std_logic;
signal heap_bh30_w3_4 :  std_logic;
signal heap_bh30_w4_4 :  std_logic;
signal CompressorIn_bh30_18_36 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_18_37 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_18_18 :  std_logic_vector(2 downto 0);
signal heap_bh30_w6_7 :  std_logic;
signal heap_bh30_w7_6 :  std_logic;
signal heap_bh30_w8_7 :  std_logic;
signal CompressorIn_bh30_19_38 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_19_39 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_19_19 :  std_logic_vector(2 downto 0);
signal heap_bh30_w9_7 :  std_logic;
signal heap_bh30_w10_6 :  std_logic;
signal heap_bh30_w11_7 :  std_logic;
signal CompressorIn_bh30_20_40 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_20_41 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_20_20 :  std_logic_vector(2 downto 0);
signal heap_bh30_w12_7 :  std_logic;
signal heap_bh30_w13_7 :  std_logic;
signal heap_bh30_w14_8 :  std_logic;
signal CompressorIn_bh30_21_42 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_21_43 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_21_21 :  std_logic_vector(2 downto 0);
signal heap_bh30_w15_8 :  std_logic;
signal heap_bh30_w16_7 :  std_logic;
signal heap_bh30_w17_8 :  std_logic;
signal CompressorIn_bh30_22_44 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_22_45 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_22_22 :  std_logic_vector(2 downto 0);
signal heap_bh30_w18_8 :  std_logic;
signal heap_bh30_w19_7 :  std_logic;
signal heap_bh30_w20_8 :  std_logic;
signal CompressorIn_bh30_23_46 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_23_47 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_23_23 :  std_logic_vector(2 downto 0);
signal heap_bh30_w21_8 :  std_logic;
signal heap_bh30_w22_7 :  std_logic;
signal heap_bh30_w23_9 :  std_logic;
signal CompressorIn_bh30_24_48 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_24_49 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_24_24 :  std_logic_vector(2 downto 0);
signal heap_bh30_w24_9 :  std_logic;
signal heap_bh30_w25_8 :  std_logic;
signal heap_bh30_w26_9 :  std_logic;
signal CompressorIn_bh30_25_50 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_25_51 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_25_25 :  std_logic_vector(2 downto 0);
signal heap_bh30_w27_9 :  std_logic;
signal heap_bh30_w28_8 :  std_logic;
signal heap_bh30_w29_9 :  std_logic;
signal CompressorIn_bh30_26_52 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_26_53 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_26_26 :  std_logic_vector(2 downto 0);
signal heap_bh30_w30_9 :  std_logic;
signal heap_bh30_w31_8 :  std_logic;
signal heap_bh30_w32_9 :  std_logic;
signal CompressorIn_bh30_27_54 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_27_55 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_27_27 :  std_logic_vector(2 downto 0);
signal heap_bh30_w33_9 :  std_logic;
signal heap_bh30_w34_8 :  std_logic;
signal heap_bh30_w35_9 :  std_logic;
signal CompressorIn_bh30_28_56 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_28_57 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_28_28 :  std_logic_vector(2 downto 0);
signal heap_bh30_w36_9 :  std_logic;
signal heap_bh30_w37_9 :  std_logic;
signal heap_bh30_w38_10 :  std_logic;
signal CompressorIn_bh30_29_58 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_29_59 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_29_29 :  std_logic_vector(2 downto 0);
signal heap_bh30_w39_10 :  std_logic;
signal heap_bh30_w40_9 :  std_logic;
signal heap_bh30_w41_10 :  std_logic;
signal CompressorIn_bh30_30_60 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_30_61 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_30_30 :  std_logic_vector(2 downto 0);
signal heap_bh30_w42_10 :  std_logic;
signal heap_bh30_w43_9 :  std_logic;
signal heap_bh30_w44_10 :  std_logic;
signal CompressorIn_bh30_31_62 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_31_63 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_31_31 :  std_logic_vector(2 downto 0);
signal heap_bh30_w45_10 :  std_logic;
signal heap_bh30_w46_9 :  std_logic;
signal heap_bh30_w47_10 :  std_logic;
signal CompressorIn_bh30_32_64 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_32_65 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_32_32 :  std_logic_vector(2 downto 0);
signal heap_bh30_w48_10 :  std_logic;
signal heap_bh30_w49_9 :  std_logic;
signal heap_bh30_w50_10 :  std_logic;
signal CompressorIn_bh30_33_66 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_33_67 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_33_33 :  std_logic_vector(2 downto 0);
signal heap_bh30_w51_10 :  std_logic;
signal heap_bh30_w52_9 :  std_logic;
signal heap_bh30_w53_10 :  std_logic;
signal CompressorIn_bh30_34_68 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_34_69 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_34_34 :  std_logic_vector(2 downto 0);
signal heap_bh30_w54_10 :  std_logic;
signal heap_bh30_w55_9 :  std_logic;
signal heap_bh30_w56_8 :  std_logic;
signal CompressorIn_bh30_35_70 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_35_71 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_35_35 :  std_logic_vector(2 downto 0);
signal heap_bh30_w56_9 :  std_logic;
signal heap_bh30_w57_8 :  std_logic;
signal heap_bh30_w58_6 :  std_logic;
signal CompressorIn_bh30_36_72 :  std_logic_vector(2 downto 0);
signal CompressorOut_bh30_36_36 :  std_logic_vector(1 downto 0);
signal heap_bh30_w4_5 :  std_logic;
signal heap_bh30_w5_6 :  std_logic;
signal CompressorIn_bh30_37_73 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_37_74 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_37_37 :  std_logic_vector(2 downto 0);
signal heap_bh30_w7_7 :  std_logic;
signal heap_bh30_w8_8 :  std_logic;
signal heap_bh30_w9_8 :  std_logic;
signal CompressorIn_bh30_38_75 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_38_76 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_38_38 :  std_logic_vector(2 downto 0);
signal heap_bh30_w10_7 :  std_logic;
signal heap_bh30_w11_8 :  std_logic;
signal heap_bh30_w12_8 :  std_logic;
signal CompressorIn_bh30_39_77 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_39_78 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_39_39 :  std_logic_vector(2 downto 0);
signal heap_bh30_w13_8 :  std_logic;
signal heap_bh30_w14_9 :  std_logic;
signal heap_bh30_w15_9 :  std_logic;
signal CompressorIn_bh30_40_79 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_40_80 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_40_40 :  std_logic_vector(2 downto 0);
signal heap_bh30_w16_8 :  std_logic;
signal heap_bh30_w17_9 :  std_logic;
signal heap_bh30_w18_9 :  std_logic;
signal CompressorIn_bh30_41_81 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_41_82 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_41_41 :  std_logic_vector(2 downto 0);
signal heap_bh30_w19_8 :  std_logic;
signal heap_bh30_w20_9 :  std_logic;
signal heap_bh30_w21_9 :  std_logic;
signal CompressorIn_bh30_42_83 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_42_84 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_42_42 :  std_logic_vector(2 downto 0);
signal heap_bh30_w22_8 :  std_logic;
signal heap_bh30_w23_10 :  std_logic;
signal heap_bh30_w24_10 :  std_logic;
signal CompressorIn_bh30_43_85 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_43_86 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_43_43 :  std_logic_vector(2 downto 0);
signal heap_bh30_w25_9 :  std_logic;
signal heap_bh30_w26_10 :  std_logic;
signal heap_bh30_w27_10 :  std_logic;
signal CompressorIn_bh30_44_87 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_44_88 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_44_44 :  std_logic_vector(2 downto 0);
signal heap_bh30_w28_9 :  std_logic;
signal heap_bh30_w29_10 :  std_logic;
signal heap_bh30_w30_10 :  std_logic;
signal CompressorIn_bh30_45_89 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_45_90 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_45_45 :  std_logic_vector(2 downto 0);
signal heap_bh30_w31_9 :  std_logic;
signal heap_bh30_w32_10 :  std_logic;
signal heap_bh30_w33_10 :  std_logic;
signal CompressorIn_bh30_46_91 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_46_92 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_46_46 :  std_logic_vector(2 downto 0);
signal heap_bh30_w34_9 :  std_logic;
signal heap_bh30_w35_10 :  std_logic;
signal heap_bh30_w36_10 :  std_logic;
signal CompressorIn_bh30_47_93 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_47_94 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_47_47 :  std_logic_vector(2 downto 0);
signal heap_bh30_w37_10 :  std_logic;
signal heap_bh30_w38_11 :  std_logic;
signal heap_bh30_w39_11 :  std_logic;
signal CompressorIn_bh30_48_95 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_48_96 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_48_48 :  std_logic_vector(2 downto 0);
signal heap_bh30_w40_10 :  std_logic;
signal heap_bh30_w41_11 :  std_logic;
signal heap_bh30_w42_11 :  std_logic;
signal CompressorIn_bh30_49_97 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_49_98 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_49_49 :  std_logic_vector(2 downto 0);
signal heap_bh30_w43_10 :  std_logic;
signal heap_bh30_w44_11 :  std_logic;
signal heap_bh30_w45_11 :  std_logic;
signal CompressorIn_bh30_50_99 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_50_100 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_50_50 :  std_logic_vector(2 downto 0);
signal heap_bh30_w46_10 :  std_logic;
signal heap_bh30_w47_11 :  std_logic;
signal heap_bh30_w48_11 :  std_logic;
signal CompressorIn_bh30_51_101 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_51_102 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_51_51 :  std_logic_vector(2 downto 0);
signal heap_bh30_w49_10 :  std_logic;
signal heap_bh30_w50_11 :  std_logic;
signal heap_bh30_w51_11 :  std_logic;
signal CompressorIn_bh30_52_103 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_52_104 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_52_52 :  std_logic_vector(2 downto 0);
signal heap_bh30_w52_10 :  std_logic;
signal heap_bh30_w53_11 :  std_logic;
signal heap_bh30_w54_11 :  std_logic;
signal CompressorIn_bh30_53_105 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_53_106 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_53_53 :  std_logic_vector(2 downto 0);
signal heap_bh30_w55_10 :  std_logic;
signal heap_bh30_w56_10 :  std_logic;
signal heap_bh30_w57_9 :  std_logic;
signal CompressorIn_bh30_54_107 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_54_108 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_54_54 :  std_logic_vector(2 downto 0);
signal heap_bh30_w57_10 :  std_logic;
signal heap_bh30_w58_7 :  std_logic;
signal heap_bh30_w59_6 :  std_logic;
signal CompressorIn_bh30_55_109 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_55_110 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_55_55 :  std_logic_vector(2 downto 0);
signal heap_bh30_w9_9 :  std_logic;
signal heap_bh30_w10_8 :  std_logic;
signal heap_bh30_w11_9 :  std_logic;
signal CompressorIn_bh30_56_111 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_56_112 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_56_56 :  std_logic_vector(2 downto 0);
signal heap_bh30_w12_9 :  std_logic;
signal heap_bh30_w13_9 :  std_logic;
signal heap_bh30_w14_10 :  std_logic;
signal CompressorIn_bh30_57_113 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_57_114 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_57_57 :  std_logic_vector(2 downto 0);
signal heap_bh30_w15_10 :  std_logic;
signal heap_bh30_w16_9 :  std_logic;
signal heap_bh30_w17_10 :  std_logic;
signal CompressorIn_bh30_58_115 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_58_116 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_58_58 :  std_logic_vector(2 downto 0);
signal heap_bh30_w18_10 :  std_logic;
signal heap_bh30_w19_9 :  std_logic;
signal heap_bh30_w20_10 :  std_logic;
signal CompressorIn_bh30_59_117 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_59_118 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_59_59 :  std_logic_vector(2 downto 0);
signal heap_bh30_w21_10 :  std_logic;
signal heap_bh30_w22_9 :  std_logic;
signal heap_bh30_w23_11 :  std_logic;
signal CompressorIn_bh30_60_119 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_60_120 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_60_60 :  std_logic_vector(2 downto 0);
signal heap_bh30_w24_11 :  std_logic;
signal heap_bh30_w25_10 :  std_logic;
signal heap_bh30_w26_11 :  std_logic;
signal CompressorIn_bh30_61_121 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_61_122 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_61_61 :  std_logic_vector(2 downto 0);
signal heap_bh30_w27_11 :  std_logic;
signal heap_bh30_w28_10 :  std_logic;
signal heap_bh30_w29_11 :  std_logic;
signal CompressorIn_bh30_62_123 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_62_124 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_62_62 :  std_logic_vector(2 downto 0);
signal heap_bh30_w30_11 :  std_logic;
signal heap_bh30_w31_10 :  std_logic;
signal heap_bh30_w32_11 :  std_logic;
signal CompressorIn_bh30_63_125 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_63_126 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_63_63 :  std_logic_vector(2 downto 0);
signal heap_bh30_w33_11 :  std_logic;
signal heap_bh30_w34_10 :  std_logic;
signal heap_bh30_w35_11 :  std_logic;
signal CompressorIn_bh30_64_127 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_64_128 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_64_64 :  std_logic_vector(2 downto 0);
signal heap_bh30_w36_11 :  std_logic;
signal heap_bh30_w37_11 :  std_logic;
signal heap_bh30_w38_12 :  std_logic;
signal CompressorIn_bh30_65_129 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_65_130 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_65_65 :  std_logic_vector(2 downto 0);
signal heap_bh30_w39_12 :  std_logic;
signal heap_bh30_w40_11 :  std_logic;
signal heap_bh30_w41_12 :  std_logic;
signal CompressorIn_bh30_66_131 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_66_132 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_66_66 :  std_logic_vector(2 downto 0);
signal heap_bh30_w42_12 :  std_logic;
signal heap_bh30_w43_11 :  std_logic;
signal heap_bh30_w44_12 :  std_logic;
signal CompressorIn_bh30_67_133 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_67_134 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_67_67 :  std_logic_vector(2 downto 0);
signal heap_bh30_w45_12 :  std_logic;
signal heap_bh30_w46_11 :  std_logic;
signal heap_bh30_w47_12 :  std_logic;
signal CompressorIn_bh30_68_135 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_68_136 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_68_68 :  std_logic_vector(2 downto 0);
signal heap_bh30_w48_12 :  std_logic;
signal heap_bh30_w49_11 :  std_logic;
signal heap_bh30_w50_12 :  std_logic;
signal CompressorIn_bh30_69_137 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_69_138 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_69_69 :  std_logic_vector(2 downto 0);
signal heap_bh30_w51_12 :  std_logic;
signal heap_bh30_w52_11 :  std_logic;
signal heap_bh30_w53_12 :  std_logic;
signal CompressorIn_bh30_70_139 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_70_140 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_70_70 :  std_logic_vector(2 downto 0);
signal heap_bh30_w54_12 :  std_logic;
signal heap_bh30_w55_11 :  std_logic;
signal heap_bh30_w56_11 :  std_logic;
signal CompressorIn_bh30_71_141 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_71_71 :  std_logic_vector(2 downto 0);
signal heap_bh30_w23_12 :  std_logic;
signal heap_bh30_w24_12 :  std_logic;
signal heap_bh30_w25_11 :  std_logic;
signal CompressorIn_bh30_72_142 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_72_72 :  std_logic_vector(2 downto 0);
signal heap_bh30_w26_12 :  std_logic;
signal heap_bh30_w27_12 :  std_logic;
signal heap_bh30_w28_11 :  std_logic;
signal CompressorIn_bh30_73_143 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_73_73 :  std_logic_vector(2 downto 0);
signal heap_bh30_w29_12 :  std_logic;
signal heap_bh30_w30_12 :  std_logic;
signal heap_bh30_w31_11 :  std_logic;
signal CompressorIn_bh30_74_144 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_74_74 :  std_logic_vector(2 downto 0);
signal heap_bh30_w32_12 :  std_logic;
signal heap_bh30_w33_12 :  std_logic;
signal heap_bh30_w34_11 :  std_logic;
signal CompressorIn_bh30_75_145 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_75_75 :  std_logic_vector(2 downto 0);
signal heap_bh30_w35_12 :  std_logic;
signal heap_bh30_w36_12 :  std_logic;
signal heap_bh30_w37_12 :  std_logic;
signal CompressorIn_bh30_76_146 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_76_76 :  std_logic_vector(2 downto 0);
signal heap_bh30_w37_13 :  std_logic;
signal heap_bh30_w38_13 :  std_logic;
signal heap_bh30_w39_13 :  std_logic;
signal CompressorIn_bh30_77_147 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_77_77 :  std_logic_vector(2 downto 0);
signal heap_bh30_w38_14 :  std_logic;
signal heap_bh30_w39_14 :  std_logic;
signal heap_bh30_w40_12 :  std_logic;
signal CompressorIn_bh30_78_148 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_78_78 :  std_logic_vector(2 downto 0);
signal heap_bh30_w39_15 :  std_logic;
signal heap_bh30_w40_13 :  std_logic;
signal heap_bh30_w41_13 :  std_logic;
signal CompressorIn_bh30_79_149 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_79_79 :  std_logic_vector(2 downto 0);
signal heap_bh30_w40_14 :  std_logic;
signal heap_bh30_w41_14 :  std_logic;
signal heap_bh30_w42_13 :  std_logic;
signal CompressorIn_bh30_80_150 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_80_80 :  std_logic_vector(2 downto 0);
signal heap_bh30_w41_15 :  std_logic;
signal heap_bh30_w42_14 :  std_logic;
signal heap_bh30_w43_12 :  std_logic;
signal CompressorIn_bh30_81_151 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_81_81 :  std_logic_vector(2 downto 0);
signal heap_bh30_w42_15 :  std_logic;
signal heap_bh30_w43_13 :  std_logic;
signal heap_bh30_w44_13 :  std_logic;
signal CompressorIn_bh30_82_152 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_82_82 :  std_logic_vector(2 downto 0);
signal heap_bh30_w43_14 :  std_logic;
signal heap_bh30_w44_14 :  std_logic;
signal heap_bh30_w45_13 :  std_logic;
signal CompressorIn_bh30_83_153 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_83_83 :  std_logic_vector(2 downto 0);
signal heap_bh30_w44_15 :  std_logic;
signal heap_bh30_w45_14 :  std_logic;
signal heap_bh30_w46_12 :  std_logic;
signal CompressorIn_bh30_84_154 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_84_84 :  std_logic_vector(2 downto 0);
signal heap_bh30_w45_15 :  std_logic;
signal heap_bh30_w46_13 :  std_logic;
signal heap_bh30_w47_13 :  std_logic;
signal CompressorIn_bh30_85_155 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_85_85 :  std_logic_vector(2 downto 0);
signal heap_bh30_w46_14 :  std_logic;
signal heap_bh30_w47_14 :  std_logic;
signal heap_bh30_w48_13 :  std_logic;
signal CompressorIn_bh30_86_156 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_86_86 :  std_logic_vector(2 downto 0);
signal heap_bh30_w47_15 :  std_logic;
signal heap_bh30_w48_14 :  std_logic;
signal heap_bh30_w49_12 :  std_logic;
signal CompressorIn_bh30_87_157 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_87_87 :  std_logic_vector(2 downto 0);
signal heap_bh30_w48_15 :  std_logic;
signal heap_bh30_w49_13 :  std_logic;
signal heap_bh30_w50_13 :  std_logic;
signal CompressorIn_bh30_88_158 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_88_88 :  std_logic_vector(2 downto 0);
signal heap_bh30_w49_14 :  std_logic;
signal heap_bh30_w50_14 :  std_logic;
signal heap_bh30_w51_13 :  std_logic;
signal CompressorIn_bh30_89_159 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_89_89 :  std_logic_vector(2 downto 0);
signal heap_bh30_w50_15 :  std_logic;
signal heap_bh30_w51_14 :  std_logic;
signal heap_bh30_w52_12 :  std_logic;
signal CompressorIn_bh30_90_160 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_90_90 :  std_logic_vector(2 downto 0);
signal heap_bh30_w51_15 :  std_logic;
signal heap_bh30_w52_13 :  std_logic;
signal heap_bh30_w53_13 :  std_logic;
signal CompressorIn_bh30_91_161 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_91_91 :  std_logic_vector(2 downto 0);
signal heap_bh30_w52_14 :  std_logic;
signal heap_bh30_w53_14 :  std_logic;
signal heap_bh30_w54_13 :  std_logic;
signal CompressorIn_bh30_92_162 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_92_92 :  std_logic_vector(2 downto 0);
signal heap_bh30_w53_15 :  std_logic;
signal heap_bh30_w54_14 :  std_logic;
signal heap_bh30_w55_12 :  std_logic;
signal CompressorIn_bh30_93_163 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_93_93 :  std_logic_vector(2 downto 0);
signal heap_bh30_w54_15 :  std_logic;
signal heap_bh30_w55_13 :  std_logic;
signal heap_bh30_w56_12 :  std_logic;
signal CompressorIn_bh30_94_164 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_94_94 :  std_logic_vector(2 downto 0);
signal heap_bh30_w55_14 :  std_logic;
signal heap_bh30_w56_13 :  std_logic;
signal heap_bh30_w57_11 :  std_logic;
signal CompressorIn_bh30_95_165 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_95_95 :  std_logic_vector(2 downto 0);
signal heap_bh30_w56_14 :  std_logic;
signal heap_bh30_w57_12 :  std_logic;
signal heap_bh30_w58_8 :  std_logic;
signal CompressorIn_bh30_96_166 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_96_96 :  std_logic_vector(2 downto 0);
signal heap_bh30_w57_13 :  std_logic;
signal heap_bh30_w58_9 :  std_logic;
signal heap_bh30_w59_7 :  std_logic;
signal CompressorIn_bh30_97_167 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_97_97 :  std_logic_vector(2 downto 0);
signal heap_bh30_w58_10 :  std_logic;
signal heap_bh30_w59_8 :  std_logic;
signal heap_bh30_w60_6 :  std_logic;
signal CompressorIn_bh30_98_168 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_98_98 :  std_logic_vector(2 downto 0);
signal heap_bh30_w59_9 :  std_logic;
signal heap_bh30_w60_7 :  std_logic;
signal heap_bh30_w61_5 :  std_logic;
signal CompressorIn_bh30_99_169 :  std_logic_vector(5 downto 0);
signal CompressorOut_bh30_99_99 :  std_logic_vector(2 downto 0);
signal heap_bh30_w60_8 :  std_logic;
signal heap_bh30_w61_6 :  std_logic;
signal heap_bh30_w62_5 :  std_logic;
signal CompressorIn_bh30_100_170 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_100_171 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_100_100 :  std_logic_vector(2 downto 0);
signal heap_bh30_w6_8 :  std_logic;
signal heap_bh30_w7_8 :  std_logic;
signal heap_bh30_w8_9 :  std_logic;
signal CompressorIn_bh30_101_172 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_101_173 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_101_101 :  std_logic_vector(2 downto 0);
signal heap_bh30_w11_10 :  std_logic;
signal heap_bh30_w12_10 :  std_logic;
signal heap_bh30_w13_10 :  std_logic;
signal CompressorIn_bh30_102_174 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_102_175 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_102_102 :  std_logic_vector(2 downto 0);
signal heap_bh30_w13_11 :  std_logic;
signal heap_bh30_w14_11 :  std_logic;
signal heap_bh30_w15_11 :  std_logic;
signal CompressorIn_bh30_103_176 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_103_177 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_103_103 :  std_logic_vector(2 downto 0);
signal heap_bh30_w14_12 :  std_logic;
signal heap_bh30_w15_12 :  std_logic;
signal heap_bh30_w16_10 :  std_logic;
signal CompressorIn_bh30_104_178 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_104_179 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_104_104 :  std_logic_vector(2 downto 0);
signal heap_bh30_w16_11 :  std_logic;
signal heap_bh30_w17_11 :  std_logic;
signal heap_bh30_w18_11 :  std_logic;
signal CompressorIn_bh30_105_180 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_105_181 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_105_105 :  std_logic_vector(2 downto 0);
signal heap_bh30_w17_12 :  std_logic;
signal heap_bh30_w18_12 :  std_logic;
signal heap_bh30_w19_10 :  std_logic;
signal CompressorIn_bh30_106_182 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_106_183 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_106_106 :  std_logic_vector(2 downto 0);
signal heap_bh30_w19_11 :  std_logic;
signal heap_bh30_w20_11 :  std_logic;
signal heap_bh30_w21_11 :  std_logic;
signal CompressorIn_bh30_107_184 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_107_185 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_107_107 :  std_logic_vector(2 downto 0);
signal heap_bh30_w20_12 :  std_logic;
signal heap_bh30_w21_12 :  std_logic;
signal heap_bh30_w22_10 :  std_logic;
signal CompressorIn_bh30_108_186 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_108_187 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_108_108 :  std_logic_vector(2 downto 0);
signal heap_bh30_w24_13 :  std_logic;
signal heap_bh30_w25_12 :  std_logic;
signal heap_bh30_w26_13 :  std_logic;
signal CompressorIn_bh30_109_188 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_109_189 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_109_109 :  std_logic_vector(2 downto 0);
signal heap_bh30_w27_13 :  std_logic;
signal heap_bh30_w28_12 :  std_logic;
signal heap_bh30_w29_13 :  std_logic;
signal CompressorIn_bh30_110_190 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_110_191 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_110_110 :  std_logic_vector(2 downto 0);
signal heap_bh30_w30_13 :  std_logic;
signal heap_bh30_w31_12 :  std_logic;
signal heap_bh30_w32_13 :  std_logic;
signal CompressorIn_bh30_111_192 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_111_193 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_111_111 :  std_logic_vector(2 downto 0);
signal heap_bh30_w33_13 :  std_logic;
signal heap_bh30_w34_12 :  std_logic;
signal heap_bh30_w35_13 :  std_logic;
signal CompressorIn_bh30_112_194 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_112_195 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_112_112 :  std_logic_vector(2 downto 0);
signal heap_bh30_w61_7 :  std_logic;
signal heap_bh30_w62_6 :  std_logic;
signal heap_bh30_w63_5 :  std_logic;
signal CompressorIn_bh30_113_196 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_113_197 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_113_113 :  std_logic_vector(2 downto 0);
signal heap_bh30_w62_7 :  std_logic;
signal heap_bh30_w63_6 :  std_logic;
signal heap_bh30_w64_4 :  std_logic;
signal CompressorIn_bh30_114_198 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_114_199 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_114_114 :  std_logic_vector(2 downto 0);
signal heap_bh30_w63_7 :  std_logic;
signal heap_bh30_w64_5 :  std_logic;
signal heap_bh30_w65_4 :  std_logic;
signal CompressorIn_bh30_115_200 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_115_201 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_115_115 :  std_logic_vector(2 downto 0);
signal heap_bh30_w65_5 :  std_logic;
signal heap_bh30_w66_4 :  std_logic;
signal heap_bh30_w67_4 :  std_logic;
signal CompressorIn_bh30_116_202 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_116_203 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_116_116 :  std_logic_vector(2 downto 0);
signal heap_bh30_w67_5 :  std_logic;
signal heap_bh30_w68_4 :  std_logic;
signal heap_bh30_w69_4 :  std_logic;
signal CompressorIn_bh30_117_204 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_117_205 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_117_117 :  std_logic_vector(2 downto 0);
signal heap_bh30_w69_5 :  std_logic;
signal heap_bh30_w70_4 :  std_logic;
signal heap_bh30_w71_4 :  std_logic;
signal CompressorIn_bh30_118_206 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_118_207 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_118_118 :  std_logic_vector(2 downto 0);
signal heap_bh30_w71_5 :  std_logic;
signal heap_bh30_w72_4 :  std_logic;
signal heap_bh30_w73_4 :  std_logic;
signal CompressorIn_bh30_119_208 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_119_209 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_119_119 :  std_logic_vector(2 downto 0);
signal heap_bh30_w73_5 :  std_logic;
signal heap_bh30_w74_4 :  std_logic;
signal heap_bh30_w75_4 :  std_logic;
signal CompressorIn_bh30_120_210 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_120_211 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_120_120 :  std_logic_vector(2 downto 0);
signal heap_bh30_w75_5 :  std_logic;
signal heap_bh30_w76_4 :  std_logic;
signal heap_bh30_w77_4 :  std_logic;
signal CompressorIn_bh30_121_212 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_121_213 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_121_121 :  std_logic_vector(2 downto 0);
signal heap_bh30_w77_5 :  std_logic;
signal heap_bh30_w78_3 :  std_logic;
signal heap_bh30_w79_3 :  std_logic;
signal CompressorIn_bh30_122_214 :  std_logic_vector(4 downto 0);
signal CompressorOut_bh30_122_122 :  std_logic_vector(2 downto 0);
signal heap_bh30_w36_13 :  std_logic;
signal heap_bh30_w37_14 :  std_logic;
signal heap_bh30_w38_15 :  std_logic;
signal CompressorIn_bh30_123_215 :  std_logic_vector(3 downto 0);
signal CompressorOut_bh30_123_123 :  std_logic_vector(2 downto 0);
signal heap_bh30_w22_11 :  std_logic;
signal heap_bh30_w23_13 :  std_logic;
signal heap_bh30_w24_14 :  std_logic;
signal CompressorIn_bh30_124_216 :  std_logic_vector(3 downto 0);
signal CompressorOut_bh30_124_124 :  std_logic_vector(2 downto 0);
signal heap_bh30_w25_13 :  std_logic;
signal heap_bh30_w26_14 :  std_logic;
signal heap_bh30_w27_14 :  std_logic;
signal CompressorIn_bh30_125_217 :  std_logic_vector(3 downto 0);
signal CompressorOut_bh30_125_125 :  std_logic_vector(2 downto 0);
signal heap_bh30_w28_13 :  std_logic;
signal heap_bh30_w29_14 :  std_logic;
signal heap_bh30_w30_14 :  std_logic;
signal CompressorIn_bh30_126_218 :  std_logic_vector(3 downto 0);
signal CompressorOut_bh30_126_126 :  std_logic_vector(2 downto 0);
signal heap_bh30_w31_13 :  std_logic;
signal heap_bh30_w32_14 :  std_logic;
signal heap_bh30_w33_14 :  std_logic;
signal CompressorIn_bh30_127_219 :  std_logic_vector(3 downto 0);
signal CompressorOut_bh30_127_127 :  std_logic_vector(2 downto 0);
signal heap_bh30_w34_13 :  std_logic;
signal heap_bh30_w35_14 :  std_logic;
signal heap_bh30_w36_14 :  std_logic;
signal CompressorIn_bh30_128_220 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_128_221 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_128_128 :  std_logic_vector(2 downto 0);
signal heap_bh30_w3_5 :  std_logic;
signal heap_bh30_w4_6 :  std_logic;
signal heap_bh30_w5_7 :  std_logic;
signal CompressorIn_bh30_129_222 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_129_223 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_129_129 :  std_logic_vector(2 downto 0);
signal heap_bh30_w8_10 :  std_logic;
signal heap_bh30_w9_10 :  std_logic;
signal heap_bh30_w10_9 :  std_logic;
signal CompressorIn_bh30_130_224 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_130_225 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_130_130 :  std_logic_vector(2 downto 0);
signal heap_bh30_w79_4 :  std_logic;
signal heap_bh30_w80_3 :  std_logic;
signal heap_bh30_w81_3 :  std_logic;
signal CompressorIn_bh30_131_226 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_131_227 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_131_131 :  std_logic_vector(2 downto 0);
signal heap_bh30_w81_4 :  std_logic;
signal heap_bh30_w82_3 :  std_logic;
signal heap_bh30_w83_3 :  std_logic;
signal CompressorIn_bh30_132_228 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_132_229 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_132_132 :  std_logic_vector(2 downto 0);
signal heap_bh30_w83_4 :  std_logic;
signal heap_bh30_w84_3 :  std_logic;
signal heap_bh30_w85_3 :  std_logic;
signal CompressorIn_bh30_133_230 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_133_231 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_133_133 :  std_logic_vector(2 downto 0);
signal heap_bh30_w85_4 :  std_logic;
signal heap_bh30_w86_3 :  std_logic;
signal heap_bh30_w87_3 :  std_logic;
signal CompressorIn_bh30_134_232 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_134_233 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_134_134 :  std_logic_vector(2 downto 0);
signal heap_bh30_w87_4 :  std_logic;
signal heap_bh30_w88_2 :  std_logic;
signal heap_bh30_w89_2 :  std_logic;
signal CompressorIn_bh30_135_234 :  std_logic_vector(2 downto 0);
signal CompressorOut_bh30_135_135 :  std_logic_vector(1 downto 0);
signal heap_bh30_w5_8 :  std_logic;
signal heap_bh30_w6_9 :  std_logic;
signal CompressorIn_bh30_136_235 :  std_logic_vector(2 downto 0);
signal CompressorOut_bh30_136_136 :  std_logic_vector(1 downto 0);
signal heap_bh30_w10_10 :  std_logic;
signal heap_bh30_w11_11 :  std_logic;
signal CompressorIn_bh30_137_236 :  std_logic_vector(2 downto 0);
signal CompressorOut_bh30_137_137 :  std_logic_vector(1 downto 0);
signal heap_bh30_w15_13 :  std_logic;
signal heap_bh30_w16_12 :  std_logic;
signal CompressorIn_bh30_138_237 :  std_logic_vector(2 downto 0);
signal CompressorOut_bh30_138_138 :  std_logic_vector(1 downto 0);
signal heap_bh30_w18_13 :  std_logic;
signal heap_bh30_w19_12 :  std_logic;
signal CompressorIn_bh30_139_238 :  std_logic_vector(2 downto 0);
signal CompressorOut_bh30_139_139 :  std_logic_vector(1 downto 0);
signal heap_bh30_w21_13 :  std_logic;
signal heap_bh30_w22_12 :  std_logic;
signal CompressorIn_bh30_140_239 :  std_logic_vector(2 downto 0);
signal CompressorOut_bh30_140_140 :  std_logic_vector(1 downto 0);
signal heap_bh30_w64_6 :  std_logic;
signal heap_bh30_w65_6 :  std_logic;
signal CompressorIn_bh30_141_240 :  std_logic_vector(2 downto 0);
signal CompressorOut_bh30_141_141 :  std_logic_vector(1 downto 0);
signal heap_bh30_w66_5 :  std_logic;
signal heap_bh30_w67_6 :  std_logic;
signal CompressorIn_bh30_142_241 :  std_logic_vector(2 downto 0);
signal CompressorOut_bh30_142_142 :  std_logic_vector(1 downto 0);
signal heap_bh30_w68_5 :  std_logic;
signal heap_bh30_w69_6 :  std_logic;
signal CompressorIn_bh30_143_242 :  std_logic_vector(2 downto 0);
signal CompressorOut_bh30_143_143 :  std_logic_vector(1 downto 0);
signal heap_bh30_w70_5 :  std_logic;
signal heap_bh30_w71_6 :  std_logic;
signal CompressorIn_bh30_144_243 :  std_logic_vector(2 downto 0);
signal CompressorOut_bh30_144_144 :  std_logic_vector(1 downto 0);
signal heap_bh30_w72_5 :  std_logic;
signal heap_bh30_w73_6 :  std_logic;
signal CompressorIn_bh30_145_244 :  std_logic_vector(2 downto 0);
signal CompressorOut_bh30_145_145 :  std_logic_vector(1 downto 0);
signal heap_bh30_w74_5 :  std_logic;
signal heap_bh30_w75_6 :  std_logic;
signal CompressorIn_bh30_146_245 :  std_logic_vector(2 downto 0);
signal CompressorOut_bh30_146_146 :  std_logic_vector(1 downto 0);
signal heap_bh30_w76_5 :  std_logic;
signal heap_bh30_w77_6 :  std_logic;
signal CompressorIn_bh30_147_246 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_147_247 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_147_147 :  std_logic_vector(2 downto 0);
signal heap_bh30_w24_15 :  std_logic;
signal heap_bh30_w25_14 :  std_logic;
signal heap_bh30_w26_15 :  std_logic;
signal CompressorIn_bh30_148_248 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_148_249 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_148_148 :  std_logic_vector(2 downto 0);
signal heap_bh30_w27_15 :  std_logic;
signal heap_bh30_w28_14 :  std_logic;
signal heap_bh30_w29_15 :  std_logic;
signal CompressorIn_bh30_149_250 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_149_251 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_149_149 :  std_logic_vector(2 downto 0);
signal heap_bh30_w30_15 :  std_logic;
signal heap_bh30_w31_14 :  std_logic;
signal heap_bh30_w32_15 :  std_logic;
signal CompressorIn_bh30_150_252 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_150_253 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_150_150 :  std_logic_vector(2 downto 0);
signal heap_bh30_w33_15 :  std_logic;
signal heap_bh30_w34_14 :  std_logic;
signal heap_bh30_w35_15 :  std_logic;
signal CompressorIn_bh30_151_254 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_151_255 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_151_151 :  std_logic_vector(2 downto 0);
signal heap_bh30_w38_16 :  std_logic;
signal heap_bh30_w39_16 :  std_logic;
signal heap_bh30_w40_15 :  std_logic;
signal CompressorIn_bh30_152_256 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_152_257 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_152_152 :  std_logic_vector(2 downto 0);
signal heap_bh30_w41_16 :  std_logic;
signal heap_bh30_w42_16 :  std_logic;
signal heap_bh30_w43_15 :  std_logic;
signal CompressorIn_bh30_153_258 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_153_259 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_153_153 :  std_logic_vector(2 downto 0);
signal heap_bh30_w44_16 :  std_logic;
signal heap_bh30_w45_16 :  std_logic;
signal heap_bh30_w46_15 :  std_logic;
signal CompressorIn_bh30_154_260 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_154_261 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_154_154 :  std_logic_vector(2 downto 0);
signal heap_bh30_w47_16 :  std_logic;
signal heap_bh30_w48_16 :  std_logic;
signal heap_bh30_w49_15 :  std_logic;
signal CompressorIn_bh30_155_262 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_155_263 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_155_155 :  std_logic_vector(2 downto 0);
signal heap_bh30_w50_16 :  std_logic;
signal heap_bh30_w51_16 :  std_logic;
signal heap_bh30_w52_15 :  std_logic;
signal CompressorIn_bh30_156_264 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_156_265 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_156_156 :  std_logic_vector(2 downto 0);
signal heap_bh30_w53_16 :  std_logic;
signal heap_bh30_w54_16 :  std_logic;
signal heap_bh30_w55_15 :  std_logic;
signal CompressorIn_bh30_157_266 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_157_267 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_157_157 :  std_logic_vector(2 downto 0);
signal heap_bh30_w56_15 :  std_logic;
signal heap_bh30_w57_14 :  std_logic;
signal heap_bh30_w58_11 :  std_logic;
signal CompressorIn_bh30_158_268 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_158_269 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_158_158 :  std_logic_vector(2 downto 0);
signal heap_bh30_w59_10 :  std_logic;
signal heap_bh30_w60_9 :  std_logic;
signal heap_bh30_w61_8 :  std_logic;
signal CompressorIn_bh30_159_270 :  std_logic_vector(3 downto 0);
signal CompressorIn_bh30_159_271 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_159_159 :  std_logic_vector(2 downto 0);
signal heap_bh30_w61_9 :  std_logic;
signal heap_bh30_w62_8 :  std_logic;
signal heap_bh30_w63_8 :  std_logic;
signal CompressorIn_bh30_160_272 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_160_273 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_160_160 :  std_logic_vector(2 downto 0);
signal heap_bh30_w7_9 :  std_logic;
signal heap_bh30_w8_11 :  std_logic;
signal heap_bh30_w9_11 :  std_logic;
signal CompressorIn_bh30_161_274 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_161_275 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_161_161 :  std_logic_vector(2 downto 0);
signal heap_bh30_w12_11 :  std_logic;
signal heap_bh30_w13_12 :  std_logic;
signal heap_bh30_w14_13 :  std_logic;
signal CompressorIn_bh30_162_276 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_162_277 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_162_162 :  std_logic_vector(2 downto 0);
signal heap_bh30_w15_14 :  std_logic;
signal heap_bh30_w16_13 :  std_logic;
signal heap_bh30_w17_13 :  std_logic;
signal CompressorIn_bh30_163_278 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_163_279 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_163_163 :  std_logic_vector(2 downto 0);
signal heap_bh30_w18_14 :  std_logic;
signal heap_bh30_w19_13 :  std_logic;
signal heap_bh30_w20_13 :  std_logic;
signal CompressorIn_bh30_164_280 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_164_281 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_164_164 :  std_logic_vector(2 downto 0);
signal heap_bh30_w21_14 :  std_logic;
signal heap_bh30_w22_13 :  std_logic;
signal heap_bh30_w23_14 :  std_logic;
signal CompressorIn_bh30_165_282 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_165_283 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_165_165 :  std_logic_vector(2 downto 0);
signal heap_bh30_w35_16 :  std_logic;
signal heap_bh30_w36_15 :  std_logic;
signal heap_bh30_w37_15 :  std_logic;
signal CompressorIn_bh30_166_284 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_166_285 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_166_166 :  std_logic_vector(2 downto 0);
signal heap_bh30_w63_9 :  std_logic;
signal heap_bh30_w64_7 :  std_logic;
signal heap_bh30_w65_7 :  std_logic;
signal CompressorIn_bh30_167_286 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_167_287 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_167_167 :  std_logic_vector(2 downto 0);
signal heap_bh30_w65_8 :  std_logic;
signal heap_bh30_w66_6 :  std_logic;
signal heap_bh30_w67_7 :  std_logic;
signal CompressorIn_bh30_168_288 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_168_289 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_168_168 :  std_logic_vector(2 downto 0);
signal heap_bh30_w67_8 :  std_logic;
signal heap_bh30_w68_6 :  std_logic;
signal heap_bh30_w69_7 :  std_logic;
signal CompressorIn_bh30_169_290 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_169_291 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_169_169 :  std_logic_vector(2 downto 0);
signal heap_bh30_w69_8 :  std_logic;
signal heap_bh30_w70_6 :  std_logic;
signal heap_bh30_w71_7 :  std_logic;
signal CompressorIn_bh30_170_292 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_170_293 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_170_170 :  std_logic_vector(2 downto 0);
signal heap_bh30_w71_8 :  std_logic;
signal heap_bh30_w72_6 :  std_logic;
signal heap_bh30_w73_7 :  std_logic;
signal CompressorIn_bh30_171_294 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_171_295 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_171_171 :  std_logic_vector(2 downto 0);
signal heap_bh30_w73_8 :  std_logic;
signal heap_bh30_w74_6 :  std_logic;
signal heap_bh30_w75_7 :  std_logic;
signal CompressorIn_bh30_172_296 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_172_297 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_172_172 :  std_logic_vector(2 downto 0);
signal heap_bh30_w75_8 :  std_logic;
signal heap_bh30_w76_6 :  std_logic;
signal heap_bh30_w77_7 :  std_logic;
signal CompressorIn_bh30_173_298 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_173_299 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_173_173 :  std_logic_vector(2 downto 0);
signal heap_bh30_w77_8 :  std_logic;
signal heap_bh30_w78_4 :  std_logic;
signal heap_bh30_w79_5 :  std_logic;
signal CompressorIn_bh30_174_300 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_174_301 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_174_174 :  std_logic_vector(2 downto 0);
signal heap_bh30_w89_3 :  std_logic;
signal heap_bh30_w90_2 :  std_logic;
signal heap_bh30_w91_2 :  std_logic;
signal CompressorIn_bh30_175_302 :  std_logic_vector(2 downto 0);
signal CompressorOut_bh30_175_175 :  std_logic_vector(1 downto 0);
signal heap_bh30_w26_16 :  std_logic;
signal heap_bh30_w27_16 :  std_logic;
signal CompressorIn_bh30_176_303 :  std_logic_vector(2 downto 0);
signal CompressorOut_bh30_176_176 :  std_logic_vector(1 downto 0);
signal heap_bh30_w29_16 :  std_logic;
signal heap_bh30_w30_16 :  std_logic;
signal CompressorIn_bh30_177_304 :  std_logic_vector(2 downto 0);
signal CompressorOut_bh30_177_177 :  std_logic_vector(1 downto 0);
signal heap_bh30_w32_16 :  std_logic;
signal heap_bh30_w33_16 :  std_logic;
signal CompressorIn_bh30_178_305 :  std_logic_vector(2 downto 0);
signal CompressorOut_bh30_178_178 :  std_logic_vector(1 downto 0);
signal heap_bh30_w37_16 :  std_logic;
signal heap_bh30_w38_17 :  std_logic;
signal CompressorIn_bh30_179_306 :  std_logic_vector(2 downto 0);
signal CompressorOut_bh30_179_179 :  std_logic_vector(1 downto 0);
signal heap_bh30_w40_16 :  std_logic;
signal heap_bh30_w41_17 :  std_logic;
signal CompressorIn_bh30_180_307 :  std_logic_vector(2 downto 0);
signal CompressorOut_bh30_180_180 :  std_logic_vector(1 downto 0);
signal heap_bh30_w43_16 :  std_logic;
signal heap_bh30_w44_17 :  std_logic;
signal CompressorIn_bh30_181_308 :  std_logic_vector(2 downto 0);
signal CompressorOut_bh30_181_181 :  std_logic_vector(1 downto 0);
signal heap_bh30_w46_16 :  std_logic;
signal heap_bh30_w47_17 :  std_logic;
signal CompressorIn_bh30_182_309 :  std_logic_vector(2 downto 0);
signal CompressorOut_bh30_182_182 :  std_logic_vector(1 downto 0);
signal heap_bh30_w49_16 :  std_logic;
signal heap_bh30_w50_17 :  std_logic;
signal CompressorIn_bh30_183_310 :  std_logic_vector(2 downto 0);
signal CompressorOut_bh30_183_183 :  std_logic_vector(1 downto 0);
signal heap_bh30_w52_16 :  std_logic;
signal heap_bh30_w53_17 :  std_logic;
signal CompressorIn_bh30_184_311 :  std_logic_vector(2 downto 0);
signal CompressorOut_bh30_184_184 :  std_logic_vector(1 downto 0);
signal heap_bh30_w55_16 :  std_logic;
signal heap_bh30_w56_16 :  std_logic;
signal CompressorIn_bh30_185_312 :  std_logic_vector(2 downto 0);
signal CompressorOut_bh30_185_185 :  std_logic_vector(1 downto 0);
signal heap_bh30_w58_12 :  std_logic;
signal heap_bh30_w59_11 :  std_logic;
signal CompressorIn_bh30_186_313 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_186_314 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_186_186 :  std_logic_vector(2 downto 0);
signal heap_bh30_w9_12 :  std_logic;
signal heap_bh30_w10_11 :  std_logic;
signal heap_bh30_w11_12 :  std_logic;
signal CompressorIn_bh30_187_315 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_187_316 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_187_187 :  std_logic_vector(2 downto 0);
signal heap_bh30_w25_15 :  std_logic;
signal heap_bh30_w26_17 :  std_logic;
signal heap_bh30_w27_17 :  std_logic;
signal CompressorIn_bh30_188_317 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_188_318 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_188_188 :  std_logic_vector(2 downto 0);
signal heap_bh30_w28_15 :  std_logic;
signal heap_bh30_w29_17 :  std_logic;
signal heap_bh30_w30_17 :  std_logic;
signal CompressorIn_bh30_189_319 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_189_320 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_189_189 :  std_logic_vector(2 downto 0);
signal heap_bh30_w31_15 :  std_logic;
signal heap_bh30_w32_17 :  std_logic;
signal heap_bh30_w33_17 :  std_logic;
signal CompressorIn_bh30_190_321 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_190_322 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_190_190 :  std_logic_vector(2 downto 0);
signal heap_bh30_w34_15 :  std_logic;
signal heap_bh30_w35_17 :  std_logic;
signal heap_bh30_w36_16 :  std_logic;
signal CompressorIn_bh30_191_323 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_191_324 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_191_191 :  std_logic_vector(2 downto 0);
signal heap_bh30_w39_17 :  std_logic;
signal heap_bh30_w40_17 :  std_logic;
signal heap_bh30_w41_18 :  std_logic;
signal CompressorIn_bh30_192_325 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_192_326 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_192_192 :  std_logic_vector(2 downto 0);
signal heap_bh30_w42_17 :  std_logic;
signal heap_bh30_w43_17 :  std_logic;
signal heap_bh30_w44_18 :  std_logic;
signal CompressorIn_bh30_193_327 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_193_328 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_193_193 :  std_logic_vector(2 downto 0);
signal heap_bh30_w45_17 :  std_logic;
signal heap_bh30_w46_17 :  std_logic;
signal heap_bh30_w47_18 :  std_logic;
signal CompressorIn_bh30_194_329 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_194_330 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_194_194 :  std_logic_vector(2 downto 0);
signal heap_bh30_w48_17 :  std_logic;
signal heap_bh30_w49_17 :  std_logic;
signal heap_bh30_w50_18 :  std_logic;
signal CompressorIn_bh30_195_331 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_195_332 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_195_195 :  std_logic_vector(2 downto 0);
signal heap_bh30_w51_17 :  std_logic;
signal heap_bh30_w52_17 :  std_logic;
signal heap_bh30_w53_18 :  std_logic;
signal CompressorIn_bh30_196_333 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_196_334 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_196_196 :  std_logic_vector(2 downto 0);
signal heap_bh30_w54_17 :  std_logic;
signal heap_bh30_w55_17 :  std_logic;
signal heap_bh30_w56_17 :  std_logic;
signal CompressorIn_bh30_197_335 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_197_336 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_197_197 :  std_logic_vector(2 downto 0);
signal heap_bh30_w57_15 :  std_logic;
signal heap_bh30_w58_13 :  std_logic;
signal heap_bh30_w59_12 :  std_logic;
signal CompressorIn_bh30_198_337 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_198_338 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_198_198 :  std_logic_vector(2 downto 0);
signal heap_bh30_w60_10 :  std_logic;
signal heap_bh30_w61_10 :  std_logic;
signal heap_bh30_w62_9 :  std_logic;
signal CompressorIn_bh30_199_339 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_199_340 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_199_199 :  std_logic_vector(2 downto 0);
signal heap_bh30_w62_10 :  std_logic;
signal heap_bh30_w63_10 :  std_logic;
signal heap_bh30_w64_8 :  std_logic;
signal CompressorIn_bh30_200_341 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_200_342 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_200_200 :  std_logic_vector(2 downto 0);
signal heap_bh30_w79_6 :  std_logic;
signal heap_bh30_w80_4 :  std_logic;
signal heap_bh30_w81_5 :  std_logic;
signal CompressorIn_bh30_201_343 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_201_344 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_201_201 :  std_logic_vector(2 downto 0);
signal heap_bh30_w91_3 :  std_logic;
signal heap_bh30_w92_2 :  std_logic;
signal heap_bh30_w93_2 :  std_logic;
signal CompressorIn_bh30_202_345 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_202_346 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_202_202 :  std_logic_vector(2 downto 0);
signal heap_bh30_w14_14 :  std_logic;
signal heap_bh30_w15_15 :  std_logic;
signal heap_bh30_w16_14 :  std_logic;
signal CompressorIn_bh30_203_347 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_203_348 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_203_203 :  std_logic_vector(2 downto 0);
signal heap_bh30_w17_14 :  std_logic;
signal heap_bh30_w18_15 :  std_logic;
signal heap_bh30_w19_14 :  std_logic;
signal CompressorIn_bh30_204_349 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_204_350 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_204_204 :  std_logic_vector(2 downto 0);
signal heap_bh30_w20_14 :  std_logic;
signal heap_bh30_w21_15 :  std_logic;
signal heap_bh30_w22_14 :  std_logic;
signal CompressorIn_bh30_205_351 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_205_352 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_205_205 :  std_logic_vector(2 downto 0);
signal heap_bh30_w23_15 :  std_logic;
signal heap_bh30_w24_16 :  std_logic;
signal heap_bh30_w25_16 :  std_logic;
signal CompressorIn_bh30_206_353 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_206_354 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_206_206 :  std_logic_vector(2 downto 0);
signal heap_bh30_w36_17 :  std_logic;
signal heap_bh30_w37_17 :  std_logic;
signal heap_bh30_w38_18 :  std_logic;
signal CompressorIn_bh30_207_355 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_207_356 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_207_207 :  std_logic_vector(2 downto 0);
signal heap_bh30_w64_9 :  std_logic;
signal heap_bh30_w65_9 :  std_logic;
signal heap_bh30_w66_7 :  std_logic;
signal CompressorIn_bh30_208_357 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_208_358 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_208_208 :  std_logic_vector(2 downto 0);
signal heap_bh30_w81_6 :  std_logic;
signal heap_bh30_w82_4 :  std_logic;
signal heap_bh30_w83_5 :  std_logic;
signal CompressorIn_bh30_209_359 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_209_360 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_209_209 :  std_logic_vector(2 downto 0);
signal heap_bh30_w93_3 :  std_logic;
signal heap_bh30_w94_2 :  std_logic;
signal heap_bh30_w95_1 :  std_logic;
signal CompressorIn_bh30_210_361 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_210_362 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_210_210 :  std_logic_vector(2 downto 0);
signal heap_bh30_w11_13 :  std_logic;
signal heap_bh30_w12_12 :  std_logic;
signal heap_bh30_w13_13 :  std_logic;
signal CompressorIn_bh30_211_363 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_211_364 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_211_211 :  std_logic_vector(2 downto 0);
signal heap_bh30_w16_15 :  std_logic;
signal heap_bh30_w17_15 :  std_logic;
signal heap_bh30_w18_16 :  std_logic;
signal CompressorIn_bh30_212_365 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_212_366 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_212_212 :  std_logic_vector(2 downto 0);
signal heap_bh30_w19_15 :  std_logic;
signal heap_bh30_w20_15 :  std_logic;
signal heap_bh30_w21_16 :  std_logic;
signal CompressorIn_bh30_213_367 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_213_368 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_213_213 :  std_logic_vector(2 downto 0);
signal heap_bh30_w22_15 :  std_logic;
signal heap_bh30_w23_16 :  std_logic;
signal heap_bh30_w24_17 :  std_logic;
signal CompressorIn_bh30_214_369 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_214_370 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_214_214 :  std_logic_vector(2 downto 0);
signal heap_bh30_w27_18 :  std_logic;
signal heap_bh30_w28_16 :  std_logic;
signal heap_bh30_w29_18 :  std_logic;
signal CompressorIn_bh30_215_371 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_215_372 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_215_215 :  std_logic_vector(2 downto 0);
signal heap_bh30_w30_18 :  std_logic;
signal heap_bh30_w31_16 :  std_logic;
signal heap_bh30_w32_18 :  std_logic;
signal CompressorIn_bh30_216_373 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_216_374 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_216_216 :  std_logic_vector(2 downto 0);
signal heap_bh30_w33_18 :  std_logic;
signal heap_bh30_w34_16 :  std_logic;
signal heap_bh30_w35_18 :  std_logic;
signal CompressorIn_bh30_217_375 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_217_376 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_217_217 :  std_logic_vector(2 downto 0);
signal heap_bh30_w41_19 :  std_logic;
signal heap_bh30_w42_18 :  std_logic;
signal heap_bh30_w43_18 :  std_logic;
signal CompressorIn_bh30_218_377 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_218_378 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_218_218 :  std_logic_vector(2 downto 0);
signal heap_bh30_w44_19 :  std_logic;
signal heap_bh30_w45_18 :  std_logic;
signal heap_bh30_w46_18 :  std_logic;
signal CompressorIn_bh30_219_379 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_219_380 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_219_219 :  std_logic_vector(2 downto 0);
signal heap_bh30_w47_19 :  std_logic;
signal heap_bh30_w48_18 :  std_logic;
signal heap_bh30_w49_18 :  std_logic;
signal CompressorIn_bh30_220_381 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_220_382 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_220_220 :  std_logic_vector(2 downto 0);
signal heap_bh30_w50_19 :  std_logic;
signal heap_bh30_w51_18 :  std_logic;
signal heap_bh30_w52_18 :  std_logic;
signal CompressorIn_bh30_221_383 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_221_384 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_221_221 :  std_logic_vector(2 downto 0);
signal heap_bh30_w53_19 :  std_logic;
signal heap_bh30_w54_18 :  std_logic;
signal heap_bh30_w55_18 :  std_logic;
signal CompressorIn_bh30_222_385 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_222_386 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_222_222 :  std_logic_vector(2 downto 0);
signal heap_bh30_w56_18 :  std_logic;
signal heap_bh30_w57_16 :  std_logic;
signal heap_bh30_w58_14 :  std_logic;
signal CompressorIn_bh30_223_387 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_223_388 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_223_223 :  std_logic_vector(2 downto 0);
signal heap_bh30_w59_13 :  std_logic;
signal heap_bh30_w60_11 :  std_logic;
signal heap_bh30_w61_11 :  std_logic;
signal CompressorIn_bh30_224_389 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_224_390 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_224_224 :  std_logic_vector(2 downto 0);
signal heap_bh30_w83_6 :  std_logic;
signal heap_bh30_w84_4 :  std_logic;
signal heap_bh30_w85_5 :  std_logic;
signal CompressorIn_bh30_225_391 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_225_392 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_225_225 :  std_logic_vector(2 downto 0);
signal heap_bh30_w38_19 :  std_logic;
signal heap_bh30_w39_18 :  std_logic;
signal heap_bh30_w40_18 :  std_logic;
signal CompressorIn_bh30_226_393 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_226_394 :  std_logic_vector(1 downto 0);
signal CompressorOut_bh30_226_226 :  std_logic_vector(2 downto 0);
signal heap_bh30_w85_6 :  std_logic;
signal heap_bh30_w86_4 :  std_logic;
signal heap_bh30_w87_5 :  std_logic;
signal CompressorIn_bh30_227_395 :  std_logic_vector(2 downto 0);
signal CompressorIn_bh30_227_396 :  std_logic_vector(0 downto 0);
signal CompressorOut_bh30_227_227 :  std_logic_vector(2 downto 0);
signal heap_bh30_w87_6 :  std_logic;
signal heap_bh30_w88_3 :  std_logic;
signal heap_bh30_w89_4 :  std_logic;
signal finalAdderIn0_bh30 :  std_logic_vector(112 downto 0);
signal finalAdderIn1_bh30 :  std_logic_vector(112 downto 0);
signal finalAdderCin_bh30 :  std_logic;
signal finalAdderOut_bh30 :  std_logic_vector(112 downto 0);
signal CompressionResult30 :  std_logic_vector(112 downto 0);
attribute rom_extract: string;
attribute rom_style: string;
attribute rom_extract of SmallMultTableP3x3r6XuYu_comb_uid103: component is "yes";
attribute rom_extract of SmallMultTableP3x3r6XuYu_comb_uid33: component is "yes";
attribute rom_extract of SmallMultTableP3x3r6XuYu_comb_uid68: component is "yes";
attribute rom_style of SmallMultTableP3x3r6XuYu_comb_uid103: component is "distributed";
attribute rom_style of SmallMultTableP3x3r6XuYu_comb_uid33: component is "distributed";
attribute rom_style of SmallMultTableP3x3r6XuYu_comb_uid68: component is "distributed";
begin
   XX_m29 <= X ;
   YY_m29 <= Y ;
   -- code generated by IntMultiplier::buildHeapLogicOnly()
   -- buildheaplogiconly called for lsbX=32 lsbY=0 msbX=56 msbY=5
   Xp_m29b31 <= XX_m29(55 downto 32) & "";
   Yp_m29b31 <= YY_m29(4 downto 0) & "0";
   x_m29b31_0 <= Xp_m29b31(2 downto 0);
   x_m29b31_1 <= Xp_m29b31(5 downto 3);
   x_m29b31_2 <= Xp_m29b31(8 downto 6);
   x_m29b31_3 <= Xp_m29b31(11 downto 9);
   x_m29b31_4 <= Xp_m29b31(14 downto 12);
   x_m29b31_5 <= Xp_m29b31(17 downto 15);
   x_m29b31_6 <= Xp_m29b31(20 downto 18);
   x_m29b31_7 <= Xp_m29b31(23 downto 21);
   y_m29b31_0 <= Yp_m29b31(2 downto 0);
   y_m29b31_1 <= Yp_m29b31(5 downto 3);
   -- Partial product row number 0
   Y0X0_31_m29 <= y_m29b31_0 & x_m29b31_0;
   PP_m29_31X0Y0_Tbl: SmallMultTableP3x3r6XuYu_comb_uid33
      port map ( X => Y0X0_31_m29,
                 Y => PP31X0Y0_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w32_0 <= PP31X0Y0_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w33_0 <= PP31X0Y0_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w34_0 <= PP31X0Y0_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w35_0 <= PP31X0Y0_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w36_0 <= PP31X0Y0_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y0X1_31_m29 <= y_m29b31_0 & x_m29b31_1;
   PP_m29_31X1Y0_Tbl: SmallMultTableP3x3r6XuYu_comb_uid33
      port map ( X => Y0X1_31_m29,
                 Y => PP31X1Y0_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w35_1 <= PP31X1Y0_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w36_1 <= PP31X1Y0_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w37_0 <= PP31X1Y0_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w38_0 <= PP31X1Y0_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w39_0 <= PP31X1Y0_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y0X2_31_m29 <= y_m29b31_0 & x_m29b31_2;
   PP_m29_31X2Y0_Tbl: SmallMultTableP3x3r6XuYu_comb_uid33
      port map ( X => Y0X2_31_m29,
                 Y => PP31X2Y0_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w38_1 <= PP31X2Y0_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w39_1 <= PP31X2Y0_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w40_0 <= PP31X2Y0_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w41_0 <= PP31X2Y0_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w42_0 <= PP31X2Y0_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y0X3_31_m29 <= y_m29b31_0 & x_m29b31_3;
   PP_m29_31X3Y0_Tbl: SmallMultTableP3x3r6XuYu_comb_uid33
      port map ( X => Y0X3_31_m29,
                 Y => PP31X3Y0_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w41_1 <= PP31X3Y0_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w42_1 <= PP31X3Y0_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w43_0 <= PP31X3Y0_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w44_0 <= PP31X3Y0_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w45_0 <= PP31X3Y0_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y0X4_31_m29 <= y_m29b31_0 & x_m29b31_4;
   PP_m29_31X4Y0_Tbl: SmallMultTableP3x3r6XuYu_comb_uid33
      port map ( X => Y0X4_31_m29,
                 Y => PP31X4Y0_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w44_1 <= PP31X4Y0_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w45_1 <= PP31X4Y0_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w46_0 <= PP31X4Y0_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w47_0 <= PP31X4Y0_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w48_0 <= PP31X4Y0_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y0X5_31_m29 <= y_m29b31_0 & x_m29b31_5;
   PP_m29_31X5Y0_Tbl: SmallMultTableP3x3r6XuYu_comb_uid33
      port map ( X => Y0X5_31_m29,
                 Y => PP31X5Y0_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w47_1 <= PP31X5Y0_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w48_1 <= PP31X5Y0_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w49_0 <= PP31X5Y0_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w50_0 <= PP31X5Y0_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w51_0 <= PP31X5Y0_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y0X6_31_m29 <= y_m29b31_0 & x_m29b31_6;
   PP_m29_31X6Y0_Tbl: SmallMultTableP3x3r6XuYu_comb_uid33
      port map ( X => Y0X6_31_m29,
                 Y => PP31X6Y0_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w50_1 <= PP31X6Y0_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w51_1 <= PP31X6Y0_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w52_0 <= PP31X6Y0_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w53_0 <= PP31X6Y0_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w54_0 <= PP31X6Y0_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y0X7_31_m29 <= y_m29b31_0 & x_m29b31_7;
   PP_m29_31X7Y0_Tbl: SmallMultTableP3x3r6XuYu_comb_uid33
      port map ( X => Y0X7_31_m29,
                 Y => PP31X7Y0_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w53_1 <= PP31X7Y0_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w54_1 <= PP31X7Y0_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w55_0 <= PP31X7Y0_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w56_0 <= PP31X7Y0_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w57_0 <= PP31X7Y0_m29(5); -- cycle= 0 cp= 5.9176e-10

   -- Partial product row number 1
   Y1X0_31_m29 <= y_m29b31_1 & x_m29b31_0;
   PP_m29_31X0Y1_Tbl: SmallMultTableP3x3r6XuYu_comb_uid33
      port map ( X => Y1X0_31_m29,
                 Y => PP31X0Y1_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w34_1 <= PP31X0Y1_m29(0); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w35_2 <= PP31X0Y1_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w36_2 <= PP31X0Y1_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w37_1 <= PP31X0Y1_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w38_2 <= PP31X0Y1_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w39_2 <= PP31X0Y1_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y1X1_31_m29 <= y_m29b31_1 & x_m29b31_1;
   PP_m29_31X1Y1_Tbl: SmallMultTableP3x3r6XuYu_comb_uid33
      port map ( X => Y1X1_31_m29,
                 Y => PP31X1Y1_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w37_2 <= PP31X1Y1_m29(0); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w38_3 <= PP31X1Y1_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w39_3 <= PP31X1Y1_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w40_1 <= PP31X1Y1_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w41_2 <= PP31X1Y1_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w42_2 <= PP31X1Y1_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y1X2_31_m29 <= y_m29b31_1 & x_m29b31_2;
   PP_m29_31X2Y1_Tbl: SmallMultTableP3x3r6XuYu_comb_uid33
      port map ( X => Y1X2_31_m29,
                 Y => PP31X2Y1_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w40_2 <= PP31X2Y1_m29(0); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w41_3 <= PP31X2Y1_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w42_3 <= PP31X2Y1_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w43_1 <= PP31X2Y1_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w44_2 <= PP31X2Y1_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w45_2 <= PP31X2Y1_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y1X3_31_m29 <= y_m29b31_1 & x_m29b31_3;
   PP_m29_31X3Y1_Tbl: SmallMultTableP3x3r6XuYu_comb_uid33
      port map ( X => Y1X3_31_m29,
                 Y => PP31X3Y1_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w43_2 <= PP31X3Y1_m29(0); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w44_3 <= PP31X3Y1_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w45_3 <= PP31X3Y1_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w46_1 <= PP31X3Y1_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w47_2 <= PP31X3Y1_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w48_2 <= PP31X3Y1_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y1X4_31_m29 <= y_m29b31_1 & x_m29b31_4;
   PP_m29_31X4Y1_Tbl: SmallMultTableP3x3r6XuYu_comb_uid33
      port map ( X => Y1X4_31_m29,
                 Y => PP31X4Y1_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w46_2 <= PP31X4Y1_m29(0); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w47_3 <= PP31X4Y1_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w48_3 <= PP31X4Y1_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w49_1 <= PP31X4Y1_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w50_2 <= PP31X4Y1_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w51_2 <= PP31X4Y1_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y1X5_31_m29 <= y_m29b31_1 & x_m29b31_5;
   PP_m29_31X5Y1_Tbl: SmallMultTableP3x3r6XuYu_comb_uid33
      port map ( X => Y1X5_31_m29,
                 Y => PP31X5Y1_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w49_2 <= PP31X5Y1_m29(0); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w50_3 <= PP31X5Y1_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w51_3 <= PP31X5Y1_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w52_1 <= PP31X5Y1_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w53_2 <= PP31X5Y1_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w54_2 <= PP31X5Y1_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y1X6_31_m29 <= y_m29b31_1 & x_m29b31_6;
   PP_m29_31X6Y1_Tbl: SmallMultTableP3x3r6XuYu_comb_uid33
      port map ( X => Y1X6_31_m29,
                 Y => PP31X6Y1_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w52_2 <= PP31X6Y1_m29(0); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w53_3 <= PP31X6Y1_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w54_3 <= PP31X6Y1_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w55_1 <= PP31X6Y1_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w56_1 <= PP31X6Y1_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w57_1 <= PP31X6Y1_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y1X7_31_m29 <= y_m29b31_1 & x_m29b31_7;
   PP_m29_31X7Y1_Tbl: SmallMultTableP3x3r6XuYu_comb_uid33
      port map ( X => Y1X7_31_m29,
                 Y => PP31X7Y1_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w55_2 <= PP31X7Y1_m29(0); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w56_2 <= PP31X7Y1_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w57_2 <= PP31X7Y1_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w58_0 <= PP31X7Y1_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w59_0 <= PP31X7Y1_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w60_0 <= PP31X7Y1_m29(5); -- cycle= 0 cp= 5.9176e-10

   -- code generated by IntMultiplier::buildHeapLogicOnly()
   -- buildheaplogiconly called for lsbX=8 lsbY=0 msbX=32 msbY=5
   Xp_m29b66 <= XX_m29(31 downto 8) & "";
   Yp_m29b66 <= YY_m29(4 downto 0) & "0";
   x_m29b66_0 <= Xp_m29b66(2 downto 0);
   x_m29b66_1 <= Xp_m29b66(5 downto 3);
   x_m29b66_2 <= Xp_m29b66(8 downto 6);
   x_m29b66_3 <= Xp_m29b66(11 downto 9);
   x_m29b66_4 <= Xp_m29b66(14 downto 12);
   x_m29b66_5 <= Xp_m29b66(17 downto 15);
   x_m29b66_6 <= Xp_m29b66(20 downto 18);
   x_m29b66_7 <= Xp_m29b66(23 downto 21);
   y_m29b66_0 <= Yp_m29b66(2 downto 0);
   y_m29b66_1 <= Yp_m29b66(5 downto 3);
   -- Partial product row number 0
   Y0X0_66_m29 <= y_m29b66_0 & x_m29b66_0;
   PP_m29_66X0Y0_Tbl: SmallMultTableP3x3r6XuYu_comb_uid68
      port map ( X => Y0X0_66_m29,
                 Y => PP66X0Y0_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w8_0 <= PP66X0Y0_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w9_0 <= PP66X0Y0_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w10_0 <= PP66X0Y0_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w11_0 <= PP66X0Y0_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w12_0 <= PP66X0Y0_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y0X1_66_m29 <= y_m29b66_0 & x_m29b66_1;
   PP_m29_66X1Y0_Tbl: SmallMultTableP3x3r6XuYu_comb_uid68
      port map ( X => Y0X1_66_m29,
                 Y => PP66X1Y0_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w11_1 <= PP66X1Y0_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w12_1 <= PP66X1Y0_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w13_0 <= PP66X1Y0_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w14_0 <= PP66X1Y0_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w15_0 <= PP66X1Y0_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y0X2_66_m29 <= y_m29b66_0 & x_m29b66_2;
   PP_m29_66X2Y0_Tbl: SmallMultTableP3x3r6XuYu_comb_uid68
      port map ( X => Y0X2_66_m29,
                 Y => PP66X2Y0_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w14_1 <= PP66X2Y0_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w15_1 <= PP66X2Y0_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w16_0 <= PP66X2Y0_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w17_0 <= PP66X2Y0_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w18_0 <= PP66X2Y0_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y0X3_66_m29 <= y_m29b66_0 & x_m29b66_3;
   PP_m29_66X3Y0_Tbl: SmallMultTableP3x3r6XuYu_comb_uid68
      port map ( X => Y0X3_66_m29,
                 Y => PP66X3Y0_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w17_1 <= PP66X3Y0_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w18_1 <= PP66X3Y0_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w19_0 <= PP66X3Y0_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w20_0 <= PP66X3Y0_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w21_0 <= PP66X3Y0_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y0X4_66_m29 <= y_m29b66_0 & x_m29b66_4;
   PP_m29_66X4Y0_Tbl: SmallMultTableP3x3r6XuYu_comb_uid68
      port map ( X => Y0X4_66_m29,
                 Y => PP66X4Y0_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w20_1 <= PP66X4Y0_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w21_1 <= PP66X4Y0_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w22_0 <= PP66X4Y0_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w23_0 <= PP66X4Y0_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w24_0 <= PP66X4Y0_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y0X5_66_m29 <= y_m29b66_0 & x_m29b66_5;
   PP_m29_66X5Y0_Tbl: SmallMultTableP3x3r6XuYu_comb_uid68
      port map ( X => Y0X5_66_m29,
                 Y => PP66X5Y0_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w23_1 <= PP66X5Y0_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w24_1 <= PP66X5Y0_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w25_0 <= PP66X5Y0_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w26_0 <= PP66X5Y0_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w27_0 <= PP66X5Y0_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y0X6_66_m29 <= y_m29b66_0 & x_m29b66_6;
   PP_m29_66X6Y0_Tbl: SmallMultTableP3x3r6XuYu_comb_uid68
      port map ( X => Y0X6_66_m29,
                 Y => PP66X6Y0_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w26_1 <= PP66X6Y0_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w27_1 <= PP66X6Y0_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w28_0 <= PP66X6Y0_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w29_0 <= PP66X6Y0_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w30_0 <= PP66X6Y0_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y0X7_66_m29 <= y_m29b66_0 & x_m29b66_7;
   PP_m29_66X7Y0_Tbl: SmallMultTableP3x3r6XuYu_comb_uid68
      port map ( X => Y0X7_66_m29,
                 Y => PP66X7Y0_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w29_1 <= PP66X7Y0_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w30_1 <= PP66X7Y0_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w31_0 <= PP66X7Y0_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w32_1 <= PP66X7Y0_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w33_1 <= PP66X7Y0_m29(5); -- cycle= 0 cp= 5.9176e-10

   -- Partial product row number 1
   Y1X0_66_m29 <= y_m29b66_1 & x_m29b66_0;
   PP_m29_66X0Y1_Tbl: SmallMultTableP3x3r6XuYu_comb_uid68
      port map ( X => Y1X0_66_m29,
                 Y => PP66X0Y1_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w10_1 <= PP66X0Y1_m29(0); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w11_2 <= PP66X0Y1_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w12_2 <= PP66X0Y1_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w13_1 <= PP66X0Y1_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w14_2 <= PP66X0Y1_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w15_2 <= PP66X0Y1_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y1X1_66_m29 <= y_m29b66_1 & x_m29b66_1;
   PP_m29_66X1Y1_Tbl: SmallMultTableP3x3r6XuYu_comb_uid68
      port map ( X => Y1X1_66_m29,
                 Y => PP66X1Y1_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w13_2 <= PP66X1Y1_m29(0); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w14_3 <= PP66X1Y1_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w15_3 <= PP66X1Y1_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w16_1 <= PP66X1Y1_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w17_2 <= PP66X1Y1_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w18_2 <= PP66X1Y1_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y1X2_66_m29 <= y_m29b66_1 & x_m29b66_2;
   PP_m29_66X2Y1_Tbl: SmallMultTableP3x3r6XuYu_comb_uid68
      port map ( X => Y1X2_66_m29,
                 Y => PP66X2Y1_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w16_2 <= PP66X2Y1_m29(0); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w17_3 <= PP66X2Y1_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w18_3 <= PP66X2Y1_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w19_1 <= PP66X2Y1_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w20_2 <= PP66X2Y1_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w21_2 <= PP66X2Y1_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y1X3_66_m29 <= y_m29b66_1 & x_m29b66_3;
   PP_m29_66X3Y1_Tbl: SmallMultTableP3x3r6XuYu_comb_uid68
      port map ( X => Y1X3_66_m29,
                 Y => PP66X3Y1_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w19_2 <= PP66X3Y1_m29(0); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w20_3 <= PP66X3Y1_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w21_3 <= PP66X3Y1_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w22_1 <= PP66X3Y1_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w23_2 <= PP66X3Y1_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w24_2 <= PP66X3Y1_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y1X4_66_m29 <= y_m29b66_1 & x_m29b66_4;
   PP_m29_66X4Y1_Tbl: SmallMultTableP3x3r6XuYu_comb_uid68
      port map ( X => Y1X4_66_m29,
                 Y => PP66X4Y1_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w22_2 <= PP66X4Y1_m29(0); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w23_3 <= PP66X4Y1_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w24_3 <= PP66X4Y1_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w25_1 <= PP66X4Y1_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w26_2 <= PP66X4Y1_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w27_2 <= PP66X4Y1_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y1X5_66_m29 <= y_m29b66_1 & x_m29b66_5;
   PP_m29_66X5Y1_Tbl: SmallMultTableP3x3r6XuYu_comb_uid68
      port map ( X => Y1X5_66_m29,
                 Y => PP66X5Y1_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w25_2 <= PP66X5Y1_m29(0); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w26_3 <= PP66X5Y1_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w27_3 <= PP66X5Y1_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w28_1 <= PP66X5Y1_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w29_2 <= PP66X5Y1_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w30_2 <= PP66X5Y1_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y1X6_66_m29 <= y_m29b66_1 & x_m29b66_6;
   PP_m29_66X6Y1_Tbl: SmallMultTableP3x3r6XuYu_comb_uid68
      port map ( X => Y1X6_66_m29,
                 Y => PP66X6Y1_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w28_2 <= PP66X6Y1_m29(0); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w29_3 <= PP66X6Y1_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w30_3 <= PP66X6Y1_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w31_1 <= PP66X6Y1_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w32_2 <= PP66X6Y1_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w33_2 <= PP66X6Y1_m29(5); -- cycle= 0 cp= 5.9176e-10

   Y1X7_66_m29 <= y_m29b66_1 & x_m29b66_7;
   PP_m29_66X7Y1_Tbl: SmallMultTableP3x3r6XuYu_comb_uid68
      port map ( X => Y1X7_66_m29,
                 Y => PP66X7Y1_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w31_2 <= PP66X7Y1_m29(0); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w32_3 <= PP66X7Y1_m29(1); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w33_3 <= PP66X7Y1_m29(2); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w34_2 <= PP66X7Y1_m29(3); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w35_3 <= PP66X7Y1_m29(4); -- cycle= 0 cp= 5.9176e-10
   heap_bh30_w36_3 <= PP66X7Y1_m29(5); -- cycle= 0 cp= 5.9176e-10

   -- code generated by IntMultiplier::buildHeapLogicOnly()
   -- buildheaplogiconly called for lsbX=0 lsbY=0 msbX=8 msbY=5
   Xp_m29b101 <= XX_m29(7 downto 0) & "0";
   Yp_m29b101 <= YY_m29(4 downto 0) & "0";
   x_m29b101_0 <= Xp_m29b101(2 downto 0);
   x_m29b101_1 <= Xp_m29b101(5 downto 3);
   x_m29b101_2 <= Xp_m29b101(8 downto 6);
   y_m29b101_0 <= Yp_m29b101(2 downto 0);
   y_m29b101_1 <= Yp_m29b101(5 downto 3);
   -- Partial product row number 0
   Y0X0_101_m29 <= y_m29b101_0 & x_m29b101_0;
   PP_m29_101X0Y0_Tbl: SmallMultTableP3x3r6XuYu_comb_uid103
      port map ( X => Y0X0_101_m29,
                 Y => PP101X0Y0_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w0_0 <= PP101X0Y0_m29(2); -- cycle= 0 cp= 5.4816e-10
   heap_bh30_w1_0 <= PP101X0Y0_m29(3); -- cycle= 0 cp= 5.4816e-10
   heap_bh30_w2_0 <= PP101X0Y0_m29(4); -- cycle= 0 cp= 5.4816e-10
   heap_bh30_w3_0 <= PP101X0Y0_m29(5); -- cycle= 0 cp= 5.4816e-10

   Y0X1_101_m29 <= y_m29b101_0 & x_m29b101_1;
   PP_m29_101X1Y0_Tbl: SmallMultTableP3x3r6XuYu_comb_uid103
      port map ( X => Y0X1_101_m29,
                 Y => PP101X1Y0_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w2_1 <= PP101X1Y0_m29(1); -- cycle= 0 cp= 5.4816e-10
   heap_bh30_w3_1 <= PP101X1Y0_m29(2); -- cycle= 0 cp= 5.4816e-10
   heap_bh30_w4_0 <= PP101X1Y0_m29(3); -- cycle= 0 cp= 5.4816e-10
   heap_bh30_w5_0 <= PP101X1Y0_m29(4); -- cycle= 0 cp= 5.4816e-10
   heap_bh30_w6_0 <= PP101X1Y0_m29(5); -- cycle= 0 cp= 5.4816e-10

   Y0X2_101_m29 <= y_m29b101_0 & x_m29b101_2;
   PP_m29_101X2Y0_Tbl: SmallMultTableP3x3r6XuYu_comb_uid103
      port map ( X => Y0X2_101_m29,
                 Y => PP101X2Y0_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w5_1 <= PP101X2Y0_m29(1); -- cycle= 0 cp= 5.4816e-10
   heap_bh30_w6_1 <= PP101X2Y0_m29(2); -- cycle= 0 cp= 5.4816e-10
   heap_bh30_w7_0 <= PP101X2Y0_m29(3); -- cycle= 0 cp= 5.4816e-10
   heap_bh30_w8_1 <= PP101X2Y0_m29(4); -- cycle= 0 cp= 5.4816e-10
   heap_bh30_w9_1 <= PP101X2Y0_m29(5); -- cycle= 0 cp= 5.4816e-10

   -- Partial product row number 1
   Y1X0_101_m29 <= y_m29b101_1 & x_m29b101_0;
   PP_m29_101X0Y1_Tbl: SmallMultTableP3x3r6XuYu_comb_uid103
      port map ( X => Y1X0_101_m29,
                 Y => PP101X0Y1_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w2_2 <= PP101X0Y1_m29(1); -- cycle= 0 cp= 5.4816e-10
   heap_bh30_w3_2 <= PP101X0Y1_m29(2); -- cycle= 0 cp= 5.4816e-10
   heap_bh30_w4_1 <= PP101X0Y1_m29(3); -- cycle= 0 cp= 5.4816e-10
   heap_bh30_w5_2 <= PP101X0Y1_m29(4); -- cycle= 0 cp= 5.4816e-10
   heap_bh30_w6_2 <= PP101X0Y1_m29(5); -- cycle= 0 cp= 5.4816e-10

   Y1X1_101_m29 <= y_m29b101_1 & x_m29b101_1;
   PP_m29_101X1Y1_Tbl: SmallMultTableP3x3r6XuYu_comb_uid103
      port map ( X => Y1X1_101_m29,
                 Y => PP101X1Y1_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w4_2 <= PP101X1Y1_m29(0); -- cycle= 0 cp= 5.4816e-10
   heap_bh30_w5_3 <= PP101X1Y1_m29(1); -- cycle= 0 cp= 5.4816e-10
   heap_bh30_w6_3 <= PP101X1Y1_m29(2); -- cycle= 0 cp= 5.4816e-10
   heap_bh30_w7_1 <= PP101X1Y1_m29(3); -- cycle= 0 cp= 5.4816e-10
   heap_bh30_w8_2 <= PP101X1Y1_m29(4); -- cycle= 0 cp= 5.4816e-10
   heap_bh30_w9_2 <= PP101X1Y1_m29(5); -- cycle= 0 cp= 5.4816e-10

   Y1X2_101_m29 <= y_m29b101_1 & x_m29b101_2;
   PP_m29_101X2Y1_Tbl: SmallMultTableP3x3r6XuYu_comb_uid103
      port map ( X => Y1X2_101_m29,
                 Y => PP101X2Y1_m29);
   -- Adding the relevant bits to the heap of bits
   heap_bh30_w7_2 <= PP101X2Y1_m29(0); -- cycle= 0 cp= 5.4816e-10
   heap_bh30_w8_3 <= PP101X2Y1_m29(1); -- cycle= 0 cp= 5.4816e-10
   heap_bh30_w9_3 <= PP101X2Y1_m29(2); -- cycle= 0 cp= 5.4816e-10
   heap_bh30_w10_2 <= PP101X2Y1_m29(3); -- cycle= 0 cp= 5.4816e-10
   heap_bh30_w11_3 <= PP101X2Y1_m29(4); -- cycle= 0 cp= 5.4816e-10
   heap_bh30_w12_3 <= PP101X2Y1_m29(5); -- cycle= 0 cp= 5.4816e-10

   
   -- Beginning of code generated by BitHeap::generateCompressorVHDL
   -- code generated by BitHeap::generateSupertileVHDL()
   DSP_bh30_ch0_0 <= std_logic_vector(unsigned("" & XX_m29(55 downto 32) & "") * unsigned("" & YY_m29(55 downto 39) & ""));
   heap_bh30_w111_0 <= DSP_bh30_ch0_0(40); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w110_0 <= DSP_bh30_ch0_0(39); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w109_0 <= DSP_bh30_ch0_0(38); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w108_0 <= DSP_bh30_ch0_0(37); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w107_0 <= DSP_bh30_ch0_0(36); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w106_0 <= DSP_bh30_ch0_0(35); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w105_0 <= DSP_bh30_ch0_0(34); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w104_0 <= DSP_bh30_ch0_0(33); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w103_0 <= DSP_bh30_ch0_0(32); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w102_0 <= DSP_bh30_ch0_0(31); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w101_0 <= DSP_bh30_ch0_0(30); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w100_0 <= DSP_bh30_ch0_0(29); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w99_0 <= DSP_bh30_ch0_0(28); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w98_0 <= DSP_bh30_ch0_0(27); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w97_0 <= DSP_bh30_ch0_0(26); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w96_0 <= DSP_bh30_ch0_0(25); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w95_0 <= DSP_bh30_ch0_0(24); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w94_0 <= DSP_bh30_ch0_0(23); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w93_0 <= DSP_bh30_ch0_0(22); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w92_0 <= DSP_bh30_ch0_0(21); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w91_0 <= DSP_bh30_ch0_0(20); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w90_0 <= DSP_bh30_ch0_0(19); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w89_0 <= DSP_bh30_ch0_0(18); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w88_0 <= DSP_bh30_ch0_0(17); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w87_0 <= DSP_bh30_ch0_0(16); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w86_0 <= DSP_bh30_ch0_0(15); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w85_0 <= DSP_bh30_ch0_0(14); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w84_0 <= DSP_bh30_ch0_0(13); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w83_0 <= DSP_bh30_ch0_0(12); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w82_0 <= DSP_bh30_ch0_0(11); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w81_0 <= DSP_bh30_ch0_0(10); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w80_0 <= DSP_bh30_ch0_0(9); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w79_0 <= DSP_bh30_ch0_0(8); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w78_0 <= DSP_bh30_ch0_0(7); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w77_0 <= DSP_bh30_ch0_0(6); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w76_0 <= DSP_bh30_ch0_0(5); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w75_0 <= DSP_bh30_ch0_0(4); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w74_0 <= DSP_bh30_ch0_0(3); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w73_0 <= DSP_bh30_ch0_0(2); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w72_0 <= DSP_bh30_ch0_0(1); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w71_0 <= DSP_bh30_ch0_0(0); -- cycle= 0 cp= 2.387e-09
   DSP_bh30_ch1_0 <= std_logic_vector(unsigned("" & XX_m29(31 downto 8) & "") * unsigned("" & YY_m29(55 downto 39) & ""));
   heap_bh30_w87_1 <= DSP_bh30_ch1_0(40); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w86_1 <= DSP_bh30_ch1_0(39); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w85_1 <= DSP_bh30_ch1_0(38); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w84_1 <= DSP_bh30_ch1_0(37); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w83_1 <= DSP_bh30_ch1_0(36); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w82_1 <= DSP_bh30_ch1_0(35); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w81_1 <= DSP_bh30_ch1_0(34); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w80_1 <= DSP_bh30_ch1_0(33); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w79_1 <= DSP_bh30_ch1_0(32); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w78_1 <= DSP_bh30_ch1_0(31); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w77_1 <= DSP_bh30_ch1_0(30); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w76_1 <= DSP_bh30_ch1_0(29); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w75_1 <= DSP_bh30_ch1_0(28); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w74_1 <= DSP_bh30_ch1_0(27); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w73_1 <= DSP_bh30_ch1_0(26); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w72_1 <= DSP_bh30_ch1_0(25); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w71_1 <= DSP_bh30_ch1_0(24); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w70_0 <= DSP_bh30_ch1_0(23); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w69_0 <= DSP_bh30_ch1_0(22); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w68_0 <= DSP_bh30_ch1_0(21); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w67_0 <= DSP_bh30_ch1_0(20); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w66_0 <= DSP_bh30_ch1_0(19); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w65_0 <= DSP_bh30_ch1_0(18); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w64_0 <= DSP_bh30_ch1_0(17); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w63_0 <= DSP_bh30_ch1_0(16); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w62_0 <= DSP_bh30_ch1_0(15); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w61_0 <= DSP_bh30_ch1_0(14); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w60_1 <= DSP_bh30_ch1_0(13); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w59_1 <= DSP_bh30_ch1_0(12); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w58_1 <= DSP_bh30_ch1_0(11); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w57_3 <= DSP_bh30_ch1_0(10); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w56_3 <= DSP_bh30_ch1_0(9); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w55_3 <= DSP_bh30_ch1_0(8); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w54_4 <= DSP_bh30_ch1_0(7); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w53_4 <= DSP_bh30_ch1_0(6); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w52_3 <= DSP_bh30_ch1_0(5); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w51_4 <= DSP_bh30_ch1_0(4); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w50_4 <= DSP_bh30_ch1_0(3); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w49_3 <= DSP_bh30_ch1_0(2); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w48_4 <= DSP_bh30_ch1_0(1); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w47_4 <= DSP_bh30_ch1_0(0); -- cycle= 0 cp= 2.387e-09
   DSP_bh30_ch2_0 <= std_logic_vector(unsigned("" & XX_m29(7 downto 0) & "0000000000000000") * unsigned("" & YY_m29(55 downto 39) & ""));
   heap_bh30_w63_1 <= DSP_bh30_ch2_0(40); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w62_1 <= DSP_bh30_ch2_0(39); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w61_1 <= DSP_bh30_ch2_0(38); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w60_2 <= DSP_bh30_ch2_0(37); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w59_2 <= DSP_bh30_ch2_0(36); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w58_2 <= DSP_bh30_ch2_0(35); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w57_4 <= DSP_bh30_ch2_0(34); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w56_4 <= DSP_bh30_ch2_0(33); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w55_4 <= DSP_bh30_ch2_0(32); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w54_5 <= DSP_bh30_ch2_0(31); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w53_5 <= DSP_bh30_ch2_0(30); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w52_4 <= DSP_bh30_ch2_0(29); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w51_5 <= DSP_bh30_ch2_0(28); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w50_5 <= DSP_bh30_ch2_0(27); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w49_4 <= DSP_bh30_ch2_0(26); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w48_5 <= DSP_bh30_ch2_0(25); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w47_5 <= DSP_bh30_ch2_0(24); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w46_3 <= DSP_bh30_ch2_0(23); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w45_4 <= DSP_bh30_ch2_0(22); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w44_4 <= DSP_bh30_ch2_0(21); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w43_3 <= DSP_bh30_ch2_0(20); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w42_4 <= DSP_bh30_ch2_0(19); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w41_4 <= DSP_bh30_ch2_0(18); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w40_3 <= DSP_bh30_ch2_0(17); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w39_4 <= DSP_bh30_ch2_0(16); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w38_4 <= DSP_bh30_ch2_0(15); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w37_3 <= DSP_bh30_ch2_0(14); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w36_4 <= DSP_bh30_ch2_0(13); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w35_4 <= DSP_bh30_ch2_0(12); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w34_3 <= DSP_bh30_ch2_0(11); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w33_4 <= DSP_bh30_ch2_0(10); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w32_4 <= DSP_bh30_ch2_0(9); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w31_3 <= DSP_bh30_ch2_0(8); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w30_4 <= DSP_bh30_ch2_0(7); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w29_4 <= DSP_bh30_ch2_0(6); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w28_3 <= DSP_bh30_ch2_0(5); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w27_4 <= DSP_bh30_ch2_0(4); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w26_4 <= DSP_bh30_ch2_0(3); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w25_3 <= DSP_bh30_ch2_0(2); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w24_4 <= DSP_bh30_ch2_0(1); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w23_4 <= DSP_bh30_ch2_0(0); -- cycle= 0 cp= 2.387e-09
   DSP_bh30_ch3_0 <= std_logic_vector(unsigned("" & XX_m29(55 downto 32) & "") * unsigned("" & YY_m29(38 downto 22) & ""));
   heap_bh30_w94_1 <= DSP_bh30_ch3_0(40); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w93_1 <= DSP_bh30_ch3_0(39); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w92_1 <= DSP_bh30_ch3_0(38); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w91_1 <= DSP_bh30_ch3_0(37); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w90_1 <= DSP_bh30_ch3_0(36); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w89_1 <= DSP_bh30_ch3_0(35); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w88_1 <= DSP_bh30_ch3_0(34); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w87_2 <= DSP_bh30_ch3_0(33); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w86_2 <= DSP_bh30_ch3_0(32); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w85_2 <= DSP_bh30_ch3_0(31); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w84_2 <= DSP_bh30_ch3_0(30); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w83_2 <= DSP_bh30_ch3_0(29); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w82_2 <= DSP_bh30_ch3_0(28); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w81_2 <= DSP_bh30_ch3_0(27); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w80_2 <= DSP_bh30_ch3_0(26); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w79_2 <= DSP_bh30_ch3_0(25); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w78_2 <= DSP_bh30_ch3_0(24); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w77_2 <= DSP_bh30_ch3_0(23); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w76_2 <= DSP_bh30_ch3_0(22); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w75_2 <= DSP_bh30_ch3_0(21); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w74_2 <= DSP_bh30_ch3_0(20); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w73_2 <= DSP_bh30_ch3_0(19); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w72_2 <= DSP_bh30_ch3_0(18); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w71_2 <= DSP_bh30_ch3_0(17); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w70_1 <= DSP_bh30_ch3_0(16); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w69_1 <= DSP_bh30_ch3_0(15); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w68_1 <= DSP_bh30_ch3_0(14); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w67_1 <= DSP_bh30_ch3_0(13); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w66_1 <= DSP_bh30_ch3_0(12); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w65_1 <= DSP_bh30_ch3_0(11); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w64_1 <= DSP_bh30_ch3_0(10); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w63_2 <= DSP_bh30_ch3_0(9); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w62_2 <= DSP_bh30_ch3_0(8); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w61_2 <= DSP_bh30_ch3_0(7); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w60_3 <= DSP_bh30_ch3_0(6); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w59_3 <= DSP_bh30_ch3_0(5); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w58_3 <= DSP_bh30_ch3_0(4); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w57_5 <= DSP_bh30_ch3_0(3); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w56_5 <= DSP_bh30_ch3_0(2); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w55_5 <= DSP_bh30_ch3_0(1); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w54_6 <= DSP_bh30_ch3_0(0); -- cycle= 0 cp= 2.387e-09
   DSP_bh30_ch4_0 <= std_logic_vector(unsigned("" & XX_m29(31 downto 8) & "") * unsigned("" & YY_m29(38 downto 22) & ""));
   heap_bh30_w70_2 <= DSP_bh30_ch4_0(40); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w69_2 <= DSP_bh30_ch4_0(39); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w68_2 <= DSP_bh30_ch4_0(38); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w67_2 <= DSP_bh30_ch4_0(37); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w66_2 <= DSP_bh30_ch4_0(36); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w65_2 <= DSP_bh30_ch4_0(35); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w64_2 <= DSP_bh30_ch4_0(34); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w63_3 <= DSP_bh30_ch4_0(33); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w62_3 <= DSP_bh30_ch4_0(32); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w61_3 <= DSP_bh30_ch4_0(31); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w60_4 <= DSP_bh30_ch4_0(30); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w59_4 <= DSP_bh30_ch4_0(29); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w58_4 <= DSP_bh30_ch4_0(28); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w57_6 <= DSP_bh30_ch4_0(27); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w56_6 <= DSP_bh30_ch4_0(26); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w55_6 <= DSP_bh30_ch4_0(25); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w54_7 <= DSP_bh30_ch4_0(24); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w53_6 <= DSP_bh30_ch4_0(23); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w52_5 <= DSP_bh30_ch4_0(22); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w51_6 <= DSP_bh30_ch4_0(21); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w50_6 <= DSP_bh30_ch4_0(20); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w49_5 <= DSP_bh30_ch4_0(19); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w48_6 <= DSP_bh30_ch4_0(18); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w47_6 <= DSP_bh30_ch4_0(17); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w46_4 <= DSP_bh30_ch4_0(16); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w45_5 <= DSP_bh30_ch4_0(15); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w44_5 <= DSP_bh30_ch4_0(14); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w43_4 <= DSP_bh30_ch4_0(13); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w42_5 <= DSP_bh30_ch4_0(12); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w41_5 <= DSP_bh30_ch4_0(11); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w40_4 <= DSP_bh30_ch4_0(10); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w39_5 <= DSP_bh30_ch4_0(9); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w38_5 <= DSP_bh30_ch4_0(8); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w37_4 <= DSP_bh30_ch4_0(7); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w36_5 <= DSP_bh30_ch4_0(6); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w35_5 <= DSP_bh30_ch4_0(5); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w34_4 <= DSP_bh30_ch4_0(4); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w33_5 <= DSP_bh30_ch4_0(3); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w32_5 <= DSP_bh30_ch4_0(2); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w31_4 <= DSP_bh30_ch4_0(1); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w30_5 <= DSP_bh30_ch4_0(0); -- cycle= 0 cp= 2.387e-09
   DSP_bh30_ch5_0 <= std_logic_vector(unsigned("" & XX_m29(7 downto 0) & "0000000000000000") * unsigned("" & YY_m29(38 downto 22) & ""));
   heap_bh30_w46_5 <= DSP_bh30_ch5_0(40); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w45_6 <= DSP_bh30_ch5_0(39); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w44_6 <= DSP_bh30_ch5_0(38); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w43_5 <= DSP_bh30_ch5_0(37); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w42_6 <= DSP_bh30_ch5_0(36); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w41_6 <= DSP_bh30_ch5_0(35); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w40_5 <= DSP_bh30_ch5_0(34); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w39_6 <= DSP_bh30_ch5_0(33); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w38_6 <= DSP_bh30_ch5_0(32); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w37_5 <= DSP_bh30_ch5_0(31); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w36_6 <= DSP_bh30_ch5_0(30); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w35_6 <= DSP_bh30_ch5_0(29); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w34_5 <= DSP_bh30_ch5_0(28); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w33_6 <= DSP_bh30_ch5_0(27); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w32_6 <= DSP_bh30_ch5_0(26); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w31_5 <= DSP_bh30_ch5_0(25); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w30_6 <= DSP_bh30_ch5_0(24); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w29_5 <= DSP_bh30_ch5_0(23); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w28_4 <= DSP_bh30_ch5_0(22); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w27_5 <= DSP_bh30_ch5_0(21); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w26_5 <= DSP_bh30_ch5_0(20); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w25_4 <= DSP_bh30_ch5_0(19); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w24_5 <= DSP_bh30_ch5_0(18); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w23_5 <= DSP_bh30_ch5_0(17); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w22_3 <= DSP_bh30_ch5_0(16); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w21_4 <= DSP_bh30_ch5_0(15); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w20_4 <= DSP_bh30_ch5_0(14); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w19_3 <= DSP_bh30_ch5_0(13); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w18_4 <= DSP_bh30_ch5_0(12); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w17_4 <= DSP_bh30_ch5_0(11); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w16_3 <= DSP_bh30_ch5_0(10); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w15_4 <= DSP_bh30_ch5_0(9); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w14_4 <= DSP_bh30_ch5_0(8); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w13_3 <= DSP_bh30_ch5_0(7); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w12_4 <= DSP_bh30_ch5_0(6); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w11_4 <= DSP_bh30_ch5_0(5); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w10_3 <= DSP_bh30_ch5_0(4); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w9_4 <= DSP_bh30_ch5_0(3); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w8_4 <= DSP_bh30_ch5_0(2); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w7_3 <= DSP_bh30_ch5_0(1); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w6_4 <= DSP_bh30_ch5_0(0); -- cycle= 0 cp= 2.387e-09
   DSP_bh30_ch6_0 <= std_logic_vector(unsigned("" & XX_m29(55 downto 32) & "") * unsigned("" & YY_m29(21 downto 5) & ""));
   heap_bh30_w77_3 <= DSP_bh30_ch6_0(40); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w76_3 <= DSP_bh30_ch6_0(39); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w75_3 <= DSP_bh30_ch6_0(38); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w74_3 <= DSP_bh30_ch6_0(37); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w73_3 <= DSP_bh30_ch6_0(36); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w72_3 <= DSP_bh30_ch6_0(35); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w71_3 <= DSP_bh30_ch6_0(34); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w70_3 <= DSP_bh30_ch6_0(33); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w69_3 <= DSP_bh30_ch6_0(32); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w68_3 <= DSP_bh30_ch6_0(31); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w67_3 <= DSP_bh30_ch6_0(30); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w66_3 <= DSP_bh30_ch6_0(29); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w65_3 <= DSP_bh30_ch6_0(28); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w64_3 <= DSP_bh30_ch6_0(27); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w63_4 <= DSP_bh30_ch6_0(26); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w62_4 <= DSP_bh30_ch6_0(25); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w61_4 <= DSP_bh30_ch6_0(24); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w60_5 <= DSP_bh30_ch6_0(23); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w59_5 <= DSP_bh30_ch6_0(22); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w58_5 <= DSP_bh30_ch6_0(21); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w57_7 <= DSP_bh30_ch6_0(20); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w56_7 <= DSP_bh30_ch6_0(19); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w55_7 <= DSP_bh30_ch6_0(18); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w54_8 <= DSP_bh30_ch6_0(17); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w53_7 <= DSP_bh30_ch6_0(16); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w52_6 <= DSP_bh30_ch6_0(15); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w51_7 <= DSP_bh30_ch6_0(14); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w50_7 <= DSP_bh30_ch6_0(13); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w49_6 <= DSP_bh30_ch6_0(12); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w48_7 <= DSP_bh30_ch6_0(11); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w47_7 <= DSP_bh30_ch6_0(10); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w46_6 <= DSP_bh30_ch6_0(9); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w45_7 <= DSP_bh30_ch6_0(8); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w44_7 <= DSP_bh30_ch6_0(7); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w43_6 <= DSP_bh30_ch6_0(6); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w42_7 <= DSP_bh30_ch6_0(5); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w41_7 <= DSP_bh30_ch6_0(4); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w40_6 <= DSP_bh30_ch6_0(3); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w39_7 <= DSP_bh30_ch6_0(2); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w38_7 <= DSP_bh30_ch6_0(1); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w37_6 <= DSP_bh30_ch6_0(0); -- cycle= 0 cp= 2.387e-09
   DSP_bh30_ch7_0 <= std_logic_vector(unsigned("" & XX_m29(31 downto 8) & "") * unsigned("" & YY_m29(21 downto 5) & ""));
   heap_bh30_w53_8 <= DSP_bh30_ch7_0(40); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w52_7 <= DSP_bh30_ch7_0(39); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w51_8 <= DSP_bh30_ch7_0(38); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w50_8 <= DSP_bh30_ch7_0(37); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w49_7 <= DSP_bh30_ch7_0(36); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w48_8 <= DSP_bh30_ch7_0(35); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w47_8 <= DSP_bh30_ch7_0(34); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w46_7 <= DSP_bh30_ch7_0(33); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w45_8 <= DSP_bh30_ch7_0(32); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w44_8 <= DSP_bh30_ch7_0(31); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w43_7 <= DSP_bh30_ch7_0(30); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w42_8 <= DSP_bh30_ch7_0(29); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w41_8 <= DSP_bh30_ch7_0(28); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w40_7 <= DSP_bh30_ch7_0(27); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w39_8 <= DSP_bh30_ch7_0(26); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w38_8 <= DSP_bh30_ch7_0(25); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w37_7 <= DSP_bh30_ch7_0(24); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w36_7 <= DSP_bh30_ch7_0(23); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w35_7 <= DSP_bh30_ch7_0(22); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w34_6 <= DSP_bh30_ch7_0(21); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w33_7 <= DSP_bh30_ch7_0(20); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w32_7 <= DSP_bh30_ch7_0(19); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w31_6 <= DSP_bh30_ch7_0(18); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w30_7 <= DSP_bh30_ch7_0(17); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w29_6 <= DSP_bh30_ch7_0(16); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w28_5 <= DSP_bh30_ch7_0(15); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w27_6 <= DSP_bh30_ch7_0(14); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w26_6 <= DSP_bh30_ch7_0(13); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w25_5 <= DSP_bh30_ch7_0(12); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w24_6 <= DSP_bh30_ch7_0(11); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w23_6 <= DSP_bh30_ch7_0(10); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w22_4 <= DSP_bh30_ch7_0(9); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w21_5 <= DSP_bh30_ch7_0(8); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w20_5 <= DSP_bh30_ch7_0(7); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w19_4 <= DSP_bh30_ch7_0(6); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w18_5 <= DSP_bh30_ch7_0(5); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w17_5 <= DSP_bh30_ch7_0(4); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w16_4 <= DSP_bh30_ch7_0(3); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w15_5 <= DSP_bh30_ch7_0(2); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w14_5 <= DSP_bh30_ch7_0(1); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w13_4 <= DSP_bh30_ch7_0(0); -- cycle= 0 cp= 2.387e-09
   DSP_bh30_ch8_0 <= std_logic_vector(unsigned("" & XX_m29(7 downto 0) & "0000000000000000") * unsigned("" & YY_m29(21 downto 5) & ""));
   heap_bh30_w29_7 <= DSP_bh30_ch8_0(40); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w28_6 <= DSP_bh30_ch8_0(39); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w27_7 <= DSP_bh30_ch8_0(38); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w26_7 <= DSP_bh30_ch8_0(37); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w25_6 <= DSP_bh30_ch8_0(36); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w24_7 <= DSP_bh30_ch8_0(35); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w23_7 <= DSP_bh30_ch8_0(34); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w22_5 <= DSP_bh30_ch8_0(33); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w21_6 <= DSP_bh30_ch8_0(32); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w20_6 <= DSP_bh30_ch8_0(31); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w19_5 <= DSP_bh30_ch8_0(30); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w18_6 <= DSP_bh30_ch8_0(29); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w17_6 <= DSP_bh30_ch8_0(28); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w16_5 <= DSP_bh30_ch8_0(27); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w15_6 <= DSP_bh30_ch8_0(26); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w14_6 <= DSP_bh30_ch8_0(25); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w13_5 <= DSP_bh30_ch8_0(24); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w12_5 <= DSP_bh30_ch8_0(23); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w11_5 <= DSP_bh30_ch8_0(22); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w10_4 <= DSP_bh30_ch8_0(21); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w9_5 <= DSP_bh30_ch8_0(20); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w8_5 <= DSP_bh30_ch8_0(19); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w7_4 <= DSP_bh30_ch8_0(18); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w6_5 <= DSP_bh30_ch8_0(17); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w5_4 <= DSP_bh30_ch8_0(16); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w4_3 <= DSP_bh30_ch8_0(15); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w3_3 <= DSP_bh30_ch8_0(14); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w2_3 <= DSP_bh30_ch8_0(13); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w1_1 <= DSP_bh30_ch8_0(12); -- cycle= 0 cp= 2.387e-09
   heap_bh30_w0_1 <= DSP_bh30_ch8_0(11); -- cycle= 0 cp= 2.387e-09

   -- Adding the constant bits
      -- All the constant bits are zero, nothing to add


   CompressorIn_bh30_0_0 <= heap_bh30_w5_3 & heap_bh30_w5_2 & heap_bh30_w5_1 & heap_bh30_w5_0;
   CompressorIn_bh30_0_1(0) <= heap_bh30_w6_3;
      Compressor_bh30_0: Compressor_14_3
      port map ( R => CompressorOut_bh30_0_0,
                 X0 => CompressorIn_bh30_0_0,
                 X1 => CompressorIn_bh30_0_1);
   heap_bh30_w5_5 <= CompressorOut_bh30_0_0(0); -- cycle= 0 cp= 1.07888e-09
   heap_bh30_w6_6 <= CompressorOut_bh30_0_0(1); -- cycle= 0 cp= 1.07888e-09
   heap_bh30_w7_5 <= CompressorOut_bh30_0_0(2); -- cycle= 0 cp= 1.07888e-09

   CompressorIn_bh30_1_2 <= heap_bh30_w8_3 & heap_bh30_w8_2 & heap_bh30_w8_1 & heap_bh30_w8_0;
   CompressorIn_bh30_1_3(0) <= heap_bh30_w9_3;
      Compressor_bh30_1: Compressor_14_3
      port map ( R => CompressorOut_bh30_1_1,
                 X0 => CompressorIn_bh30_1_2,
                 X1 => CompressorIn_bh30_1_3);
   heap_bh30_w8_6 <= CompressorOut_bh30_1_1(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w9_6 <= CompressorOut_bh30_1_1(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w10_5 <= CompressorOut_bh30_1_1(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_2_4 <= heap_bh30_w11_3 & heap_bh30_w11_2 & heap_bh30_w11_1 & heap_bh30_w11_0;
   CompressorIn_bh30_2_5(0) <= heap_bh30_w12_3;
      Compressor_bh30_2: Compressor_14_3
      port map ( R => CompressorOut_bh30_2_2,
                 X0 => CompressorIn_bh30_2_4,
                 X1 => CompressorIn_bh30_2_5);
   heap_bh30_w11_6 <= CompressorOut_bh30_2_2(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w12_6 <= CompressorOut_bh30_2_2(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w13_6 <= CompressorOut_bh30_2_2(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_3_6 <= heap_bh30_w14_3 & heap_bh30_w14_2 & heap_bh30_w14_1 & heap_bh30_w14_0;
   CompressorIn_bh30_3_7(0) <= heap_bh30_w15_3;
      Compressor_bh30_3: Compressor_14_3
      port map ( R => CompressorOut_bh30_3_3,
                 X0 => CompressorIn_bh30_3_6,
                 X1 => CompressorIn_bh30_3_7);
   heap_bh30_w14_7 <= CompressorOut_bh30_3_3(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w15_7 <= CompressorOut_bh30_3_3(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w16_6 <= CompressorOut_bh30_3_3(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_4_8 <= heap_bh30_w17_3 & heap_bh30_w17_2 & heap_bh30_w17_1 & heap_bh30_w17_0;
   CompressorIn_bh30_4_9(0) <= heap_bh30_w18_3;
      Compressor_bh30_4: Compressor_14_3
      port map ( R => CompressorOut_bh30_4_4,
                 X0 => CompressorIn_bh30_4_8,
                 X1 => CompressorIn_bh30_4_9);
   heap_bh30_w17_7 <= CompressorOut_bh30_4_4(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w18_7 <= CompressorOut_bh30_4_4(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w19_6 <= CompressorOut_bh30_4_4(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_5_10 <= heap_bh30_w20_3 & heap_bh30_w20_2 & heap_bh30_w20_1 & heap_bh30_w20_0;
   CompressorIn_bh30_5_11(0) <= heap_bh30_w21_3;
      Compressor_bh30_5: Compressor_14_3
      port map ( R => CompressorOut_bh30_5_5,
                 X0 => CompressorIn_bh30_5_10,
                 X1 => CompressorIn_bh30_5_11);
   heap_bh30_w20_7 <= CompressorOut_bh30_5_5(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w21_7 <= CompressorOut_bh30_5_5(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w22_6 <= CompressorOut_bh30_5_5(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_6_12 <= heap_bh30_w23_3 & heap_bh30_w23_2 & heap_bh30_w23_1 & heap_bh30_w23_0;
   CompressorIn_bh30_6_13(0) <= heap_bh30_w24_3;
      Compressor_bh30_6: Compressor_14_3
      port map ( R => CompressorOut_bh30_6_6,
                 X0 => CompressorIn_bh30_6_12,
                 X1 => CompressorIn_bh30_6_13);
   heap_bh30_w23_8 <= CompressorOut_bh30_6_6(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w24_8 <= CompressorOut_bh30_6_6(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w25_7 <= CompressorOut_bh30_6_6(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_7_14 <= heap_bh30_w26_3 & heap_bh30_w26_2 & heap_bh30_w26_1 & heap_bh30_w26_0;
   CompressorIn_bh30_7_15(0) <= heap_bh30_w27_3;
      Compressor_bh30_7: Compressor_14_3
      port map ( R => CompressorOut_bh30_7_7,
                 X0 => CompressorIn_bh30_7_14,
                 X1 => CompressorIn_bh30_7_15);
   heap_bh30_w26_8 <= CompressorOut_bh30_7_7(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w27_8 <= CompressorOut_bh30_7_7(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w28_7 <= CompressorOut_bh30_7_7(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_8_16 <= heap_bh30_w29_3 & heap_bh30_w29_2 & heap_bh30_w29_1 & heap_bh30_w29_0;
   CompressorIn_bh30_8_17(0) <= heap_bh30_w30_3;
      Compressor_bh30_8: Compressor_14_3
      port map ( R => CompressorOut_bh30_8_8,
                 X0 => CompressorIn_bh30_8_16,
                 X1 => CompressorIn_bh30_8_17);
   heap_bh30_w29_8 <= CompressorOut_bh30_8_8(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w30_8 <= CompressorOut_bh30_8_8(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w31_7 <= CompressorOut_bh30_8_8(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_9_18 <= heap_bh30_w32_3 & heap_bh30_w32_2 & heap_bh30_w32_1 & heap_bh30_w32_0;
   CompressorIn_bh30_9_19(0) <= heap_bh30_w33_3;
      Compressor_bh30_9: Compressor_14_3
      port map ( R => CompressorOut_bh30_9_9,
                 X0 => CompressorIn_bh30_9_18,
                 X1 => CompressorIn_bh30_9_19);
   heap_bh30_w32_8 <= CompressorOut_bh30_9_9(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w33_8 <= CompressorOut_bh30_9_9(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w34_7 <= CompressorOut_bh30_9_9(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_10_20 <= heap_bh30_w35_3 & heap_bh30_w35_2 & heap_bh30_w35_1 & heap_bh30_w35_0;
   CompressorIn_bh30_10_21(0) <= heap_bh30_w36_3;
      Compressor_bh30_10: Compressor_14_3
      port map ( R => CompressorOut_bh30_10_10,
                 X0 => CompressorIn_bh30_10_20,
                 X1 => CompressorIn_bh30_10_21);
   heap_bh30_w35_8 <= CompressorOut_bh30_10_10(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w36_8 <= CompressorOut_bh30_10_10(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w37_8 <= CompressorOut_bh30_10_10(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_11_22 <= heap_bh30_w38_3 & heap_bh30_w38_2 & heap_bh30_w38_1 & heap_bh30_w38_0;
   CompressorIn_bh30_11_23(0) <= heap_bh30_w39_3;
      Compressor_bh30_11: Compressor_14_3
      port map ( R => CompressorOut_bh30_11_11,
                 X0 => CompressorIn_bh30_11_22,
                 X1 => CompressorIn_bh30_11_23);
   heap_bh30_w38_9 <= CompressorOut_bh30_11_11(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w39_9 <= CompressorOut_bh30_11_11(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w40_8 <= CompressorOut_bh30_11_11(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_12_24 <= heap_bh30_w41_3 & heap_bh30_w41_2 & heap_bh30_w41_1 & heap_bh30_w41_0;
   CompressorIn_bh30_12_25(0) <= heap_bh30_w42_3;
      Compressor_bh30_12: Compressor_14_3
      port map ( R => CompressorOut_bh30_12_12,
                 X0 => CompressorIn_bh30_12_24,
                 X1 => CompressorIn_bh30_12_25);
   heap_bh30_w41_9 <= CompressorOut_bh30_12_12(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w42_9 <= CompressorOut_bh30_12_12(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w43_8 <= CompressorOut_bh30_12_12(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_13_26 <= heap_bh30_w44_3 & heap_bh30_w44_2 & heap_bh30_w44_1 & heap_bh30_w44_0;
   CompressorIn_bh30_13_27(0) <= heap_bh30_w45_3;
      Compressor_bh30_13: Compressor_14_3
      port map ( R => CompressorOut_bh30_13_13,
                 X0 => CompressorIn_bh30_13_26,
                 X1 => CompressorIn_bh30_13_27);
   heap_bh30_w44_9 <= CompressorOut_bh30_13_13(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w45_9 <= CompressorOut_bh30_13_13(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w46_8 <= CompressorOut_bh30_13_13(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_14_28 <= heap_bh30_w47_3 & heap_bh30_w47_2 & heap_bh30_w47_1 & heap_bh30_w47_0;
   CompressorIn_bh30_14_29(0) <= heap_bh30_w48_3;
      Compressor_bh30_14: Compressor_14_3
      port map ( R => CompressorOut_bh30_14_14,
                 X0 => CompressorIn_bh30_14_28,
                 X1 => CompressorIn_bh30_14_29);
   heap_bh30_w47_9 <= CompressorOut_bh30_14_14(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w48_9 <= CompressorOut_bh30_14_14(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w49_8 <= CompressorOut_bh30_14_14(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_15_30 <= heap_bh30_w50_3 & heap_bh30_w50_2 & heap_bh30_w50_1 & heap_bh30_w50_0;
   CompressorIn_bh30_15_31(0) <= heap_bh30_w51_3;
      Compressor_bh30_15: Compressor_14_3
      port map ( R => CompressorOut_bh30_15_15,
                 X0 => CompressorIn_bh30_15_30,
                 X1 => CompressorIn_bh30_15_31);
   heap_bh30_w50_9 <= CompressorOut_bh30_15_15(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w51_9 <= CompressorOut_bh30_15_15(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w52_8 <= CompressorOut_bh30_15_15(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_16_32 <= heap_bh30_w53_3 & heap_bh30_w53_2 & heap_bh30_w53_1 & heap_bh30_w53_0;
   CompressorIn_bh30_16_33(0) <= heap_bh30_w54_3;
      Compressor_bh30_16: Compressor_14_3
      port map ( R => CompressorOut_bh30_16_16,
                 X0 => CompressorIn_bh30_16_32,
                 X1 => CompressorIn_bh30_16_33);
   heap_bh30_w53_9 <= CompressorOut_bh30_16_16(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w54_9 <= CompressorOut_bh30_16_16(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w55_8 <= CompressorOut_bh30_16_16(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_17_34 <= heap_bh30_w2_2 & heap_bh30_w2_1 & heap_bh30_w2_0;
   CompressorIn_bh30_17_35 <= heap_bh30_w3_2 & heap_bh30_w3_1;
      Compressor_bh30_17: Compressor_23_3
      port map ( R => CompressorOut_bh30_17_17,
                 X0 => CompressorIn_bh30_17_34,
                 X1 => CompressorIn_bh30_17_35);
   heap_bh30_w2_4 <= CompressorOut_bh30_17_17(0); -- cycle= 0 cp= 1.07888e-09
   heap_bh30_w3_4 <= CompressorOut_bh30_17_17(1); -- cycle= 0 cp= 1.07888e-09
   heap_bh30_w4_4 <= CompressorOut_bh30_17_17(2); -- cycle= 0 cp= 1.07888e-09

   CompressorIn_bh30_18_36 <= heap_bh30_w6_2 & heap_bh30_w6_1 & heap_bh30_w6_0;
   CompressorIn_bh30_18_37 <= heap_bh30_w7_2 & heap_bh30_w7_1;
      Compressor_bh30_18: Compressor_23_3
      port map ( R => CompressorOut_bh30_18_18,
                 X0 => CompressorIn_bh30_18_36,
                 X1 => CompressorIn_bh30_18_37);
   heap_bh30_w6_7 <= CompressorOut_bh30_18_18(0); -- cycle= 0 cp= 1.07888e-09
   heap_bh30_w7_6 <= CompressorOut_bh30_18_18(1); -- cycle= 0 cp= 1.07888e-09
   heap_bh30_w8_7 <= CompressorOut_bh30_18_18(2); -- cycle= 0 cp= 1.07888e-09

   CompressorIn_bh30_19_38 <= heap_bh30_w9_2 & heap_bh30_w9_1 & heap_bh30_w9_0;
   CompressorIn_bh30_19_39 <= heap_bh30_w10_2 & heap_bh30_w10_1;
      Compressor_bh30_19: Compressor_23_3
      port map ( R => CompressorOut_bh30_19_19,
                 X0 => CompressorIn_bh30_19_38,
                 X1 => CompressorIn_bh30_19_39);
   heap_bh30_w9_7 <= CompressorOut_bh30_19_19(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w10_6 <= CompressorOut_bh30_19_19(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w11_7 <= CompressorOut_bh30_19_19(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_20_40 <= heap_bh30_w12_2 & heap_bh30_w12_1 & heap_bh30_w12_0;
   CompressorIn_bh30_20_41 <= heap_bh30_w13_2 & heap_bh30_w13_1;
      Compressor_bh30_20: Compressor_23_3
      port map ( R => CompressorOut_bh30_20_20,
                 X0 => CompressorIn_bh30_20_40,
                 X1 => CompressorIn_bh30_20_41);
   heap_bh30_w12_7 <= CompressorOut_bh30_20_20(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w13_7 <= CompressorOut_bh30_20_20(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w14_8 <= CompressorOut_bh30_20_20(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_21_42 <= heap_bh30_w15_2 & heap_bh30_w15_1 & heap_bh30_w15_0;
   CompressorIn_bh30_21_43 <= heap_bh30_w16_2 & heap_bh30_w16_1;
      Compressor_bh30_21: Compressor_23_3
      port map ( R => CompressorOut_bh30_21_21,
                 X0 => CompressorIn_bh30_21_42,
                 X1 => CompressorIn_bh30_21_43);
   heap_bh30_w15_8 <= CompressorOut_bh30_21_21(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w16_7 <= CompressorOut_bh30_21_21(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w17_8 <= CompressorOut_bh30_21_21(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_22_44 <= heap_bh30_w18_2 & heap_bh30_w18_1 & heap_bh30_w18_0;
   CompressorIn_bh30_22_45 <= heap_bh30_w19_2 & heap_bh30_w19_1;
      Compressor_bh30_22: Compressor_23_3
      port map ( R => CompressorOut_bh30_22_22,
                 X0 => CompressorIn_bh30_22_44,
                 X1 => CompressorIn_bh30_22_45);
   heap_bh30_w18_8 <= CompressorOut_bh30_22_22(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w19_7 <= CompressorOut_bh30_22_22(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w20_8 <= CompressorOut_bh30_22_22(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_23_46 <= heap_bh30_w21_2 & heap_bh30_w21_1 & heap_bh30_w21_0;
   CompressorIn_bh30_23_47 <= heap_bh30_w22_2 & heap_bh30_w22_1;
      Compressor_bh30_23: Compressor_23_3
      port map ( R => CompressorOut_bh30_23_23,
                 X0 => CompressorIn_bh30_23_46,
                 X1 => CompressorIn_bh30_23_47);
   heap_bh30_w21_8 <= CompressorOut_bh30_23_23(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w22_7 <= CompressorOut_bh30_23_23(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w23_9 <= CompressorOut_bh30_23_23(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_24_48 <= heap_bh30_w24_2 & heap_bh30_w24_1 & heap_bh30_w24_0;
   CompressorIn_bh30_24_49 <= heap_bh30_w25_2 & heap_bh30_w25_1;
      Compressor_bh30_24: Compressor_23_3
      port map ( R => CompressorOut_bh30_24_24,
                 X0 => CompressorIn_bh30_24_48,
                 X1 => CompressorIn_bh30_24_49);
   heap_bh30_w24_9 <= CompressorOut_bh30_24_24(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w25_8 <= CompressorOut_bh30_24_24(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w26_9 <= CompressorOut_bh30_24_24(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_25_50 <= heap_bh30_w27_2 & heap_bh30_w27_1 & heap_bh30_w27_0;
   CompressorIn_bh30_25_51 <= heap_bh30_w28_2 & heap_bh30_w28_1;
      Compressor_bh30_25: Compressor_23_3
      port map ( R => CompressorOut_bh30_25_25,
                 X0 => CompressorIn_bh30_25_50,
                 X1 => CompressorIn_bh30_25_51);
   heap_bh30_w27_9 <= CompressorOut_bh30_25_25(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w28_8 <= CompressorOut_bh30_25_25(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w29_9 <= CompressorOut_bh30_25_25(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_26_52 <= heap_bh30_w30_2 & heap_bh30_w30_1 & heap_bh30_w30_0;
   CompressorIn_bh30_26_53 <= heap_bh30_w31_2 & heap_bh30_w31_1;
      Compressor_bh30_26: Compressor_23_3
      port map ( R => CompressorOut_bh30_26_26,
                 X0 => CompressorIn_bh30_26_52,
                 X1 => CompressorIn_bh30_26_53);
   heap_bh30_w30_9 <= CompressorOut_bh30_26_26(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w31_8 <= CompressorOut_bh30_26_26(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w32_9 <= CompressorOut_bh30_26_26(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_27_54 <= heap_bh30_w33_2 & heap_bh30_w33_1 & heap_bh30_w33_0;
   CompressorIn_bh30_27_55 <= heap_bh30_w34_2 & heap_bh30_w34_1;
      Compressor_bh30_27: Compressor_23_3
      port map ( R => CompressorOut_bh30_27_27,
                 X0 => CompressorIn_bh30_27_54,
                 X1 => CompressorIn_bh30_27_55);
   heap_bh30_w33_9 <= CompressorOut_bh30_27_27(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w34_8 <= CompressorOut_bh30_27_27(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w35_9 <= CompressorOut_bh30_27_27(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_28_56 <= heap_bh30_w36_2 & heap_bh30_w36_1 & heap_bh30_w36_0;
   CompressorIn_bh30_28_57 <= heap_bh30_w37_2 & heap_bh30_w37_1;
      Compressor_bh30_28: Compressor_23_3
      port map ( R => CompressorOut_bh30_28_28,
                 X0 => CompressorIn_bh30_28_56,
                 X1 => CompressorIn_bh30_28_57);
   heap_bh30_w36_9 <= CompressorOut_bh30_28_28(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w37_9 <= CompressorOut_bh30_28_28(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w38_10 <= CompressorOut_bh30_28_28(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_29_58 <= heap_bh30_w39_2 & heap_bh30_w39_1 & heap_bh30_w39_0;
   CompressorIn_bh30_29_59 <= heap_bh30_w40_2 & heap_bh30_w40_1;
      Compressor_bh30_29: Compressor_23_3
      port map ( R => CompressorOut_bh30_29_29,
                 X0 => CompressorIn_bh30_29_58,
                 X1 => CompressorIn_bh30_29_59);
   heap_bh30_w39_10 <= CompressorOut_bh30_29_29(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w40_9 <= CompressorOut_bh30_29_29(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w41_10 <= CompressorOut_bh30_29_29(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_30_60 <= heap_bh30_w42_2 & heap_bh30_w42_1 & heap_bh30_w42_0;
   CompressorIn_bh30_30_61 <= heap_bh30_w43_2 & heap_bh30_w43_1;
      Compressor_bh30_30: Compressor_23_3
      port map ( R => CompressorOut_bh30_30_30,
                 X0 => CompressorIn_bh30_30_60,
                 X1 => CompressorIn_bh30_30_61);
   heap_bh30_w42_10 <= CompressorOut_bh30_30_30(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w43_9 <= CompressorOut_bh30_30_30(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w44_10 <= CompressorOut_bh30_30_30(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_31_62 <= heap_bh30_w45_2 & heap_bh30_w45_1 & heap_bh30_w45_0;
   CompressorIn_bh30_31_63 <= heap_bh30_w46_2 & heap_bh30_w46_1;
      Compressor_bh30_31: Compressor_23_3
      port map ( R => CompressorOut_bh30_31_31,
                 X0 => CompressorIn_bh30_31_62,
                 X1 => CompressorIn_bh30_31_63);
   heap_bh30_w45_10 <= CompressorOut_bh30_31_31(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w46_9 <= CompressorOut_bh30_31_31(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w47_10 <= CompressorOut_bh30_31_31(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_32_64 <= heap_bh30_w48_2 & heap_bh30_w48_1 & heap_bh30_w48_0;
   CompressorIn_bh30_32_65 <= heap_bh30_w49_2 & heap_bh30_w49_1;
      Compressor_bh30_32: Compressor_23_3
      port map ( R => CompressorOut_bh30_32_32,
                 X0 => CompressorIn_bh30_32_64,
                 X1 => CompressorIn_bh30_32_65);
   heap_bh30_w48_10 <= CompressorOut_bh30_32_32(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w49_9 <= CompressorOut_bh30_32_32(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w50_10 <= CompressorOut_bh30_32_32(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_33_66 <= heap_bh30_w51_2 & heap_bh30_w51_1 & heap_bh30_w51_0;
   CompressorIn_bh30_33_67 <= heap_bh30_w52_2 & heap_bh30_w52_1;
      Compressor_bh30_33: Compressor_23_3
      port map ( R => CompressorOut_bh30_33_33,
                 X0 => CompressorIn_bh30_33_66,
                 X1 => CompressorIn_bh30_33_67);
   heap_bh30_w51_10 <= CompressorOut_bh30_33_33(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w52_9 <= CompressorOut_bh30_33_33(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w53_10 <= CompressorOut_bh30_33_33(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_34_68 <= heap_bh30_w54_2 & heap_bh30_w54_1 & heap_bh30_w54_0;
   CompressorIn_bh30_34_69 <= heap_bh30_w55_2 & heap_bh30_w55_1;
      Compressor_bh30_34: Compressor_23_3
      port map ( R => CompressorOut_bh30_34_34,
                 X0 => CompressorIn_bh30_34_68,
                 X1 => CompressorIn_bh30_34_69);
   heap_bh30_w54_10 <= CompressorOut_bh30_34_34(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w55_9 <= CompressorOut_bh30_34_34(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w56_8 <= CompressorOut_bh30_34_34(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_35_70 <= heap_bh30_w56_2 & heap_bh30_w56_1 & heap_bh30_w56_0;
   CompressorIn_bh30_35_71 <= heap_bh30_w57_2 & heap_bh30_w57_1;
      Compressor_bh30_35: Compressor_23_3
      port map ( R => CompressorOut_bh30_35_35,
                 X0 => CompressorIn_bh30_35_70,
                 X1 => CompressorIn_bh30_35_71);
   heap_bh30_w56_9 <= CompressorOut_bh30_35_35(0); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w57_8 <= CompressorOut_bh30_35_35(1); -- cycle= 0 cp= 1.12248e-09
   heap_bh30_w58_6 <= CompressorOut_bh30_35_35(2); -- cycle= 0 cp= 1.12248e-09

   CompressorIn_bh30_36_72 <= heap_bh30_w4_2 & heap_bh30_w4_1 & heap_bh30_w4_0;
      Compressor_bh30_36: Compressor_3_2
      port map ( R => CompressorOut_bh30_36_36,
                 X0 => CompressorIn_bh30_36_72);
   heap_bh30_w4_5 <= CompressorOut_bh30_36_36(0); -- cycle= 0 cp= 1.07888e-09
   heap_bh30_w5_6 <= CompressorOut_bh30_36_36(1); -- cycle= 0 cp= 1.07888e-09

   CompressorIn_bh30_37_73 <= heap_bh30_w7_0 & heap_bh30_w7_6 & heap_bh30_w7_5;
   CompressorIn_bh30_37_74 <= heap_bh30_w8_7 & heap_bh30_w8_6;
      Compressor_bh30_37: Compressor_23_3
      port map ( R => CompressorOut_bh30_37_37,
                 X0 => CompressorIn_bh30_37_73,
                 X1 => CompressorIn_bh30_37_74);
   heap_bh30_w7_7 <= CompressorOut_bh30_37_37(0); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w8_8 <= CompressorOut_bh30_37_37(1); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w9_8 <= CompressorOut_bh30_37_37(2); -- cycle= 0 cp= 1.6532e-09

   CompressorIn_bh30_38_75 <= heap_bh30_w10_0 & heap_bh30_w10_6 & heap_bh30_w10_5;
   CompressorIn_bh30_38_76 <= heap_bh30_w11_7 & heap_bh30_w11_6;
      Compressor_bh30_38: Compressor_23_3
      port map ( R => CompressorOut_bh30_38_38,
                 X0 => CompressorIn_bh30_38_75,
                 X1 => CompressorIn_bh30_38_76);
   heap_bh30_w10_7 <= CompressorOut_bh30_38_38(0); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w11_8 <= CompressorOut_bh30_38_38(1); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w12_8 <= CompressorOut_bh30_38_38(2); -- cycle= 0 cp= 1.6532e-09

   CompressorIn_bh30_39_77 <= heap_bh30_w13_0 & heap_bh30_w13_7 & heap_bh30_w13_6;
   CompressorIn_bh30_39_78 <= heap_bh30_w14_8 & heap_bh30_w14_7;
      Compressor_bh30_39: Compressor_23_3
      port map ( R => CompressorOut_bh30_39_39,
                 X0 => CompressorIn_bh30_39_77,
                 X1 => CompressorIn_bh30_39_78);
   heap_bh30_w13_8 <= CompressorOut_bh30_39_39(0); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w14_9 <= CompressorOut_bh30_39_39(1); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w15_9 <= CompressorOut_bh30_39_39(2); -- cycle= 0 cp= 1.6532e-09

   CompressorIn_bh30_40_79 <= heap_bh30_w16_0 & heap_bh30_w16_7 & heap_bh30_w16_6;
   CompressorIn_bh30_40_80 <= heap_bh30_w17_8 & heap_bh30_w17_7;
      Compressor_bh30_40: Compressor_23_3
      port map ( R => CompressorOut_bh30_40_40,
                 X0 => CompressorIn_bh30_40_79,
                 X1 => CompressorIn_bh30_40_80);
   heap_bh30_w16_8 <= CompressorOut_bh30_40_40(0); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w17_9 <= CompressorOut_bh30_40_40(1); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w18_9 <= CompressorOut_bh30_40_40(2); -- cycle= 0 cp= 1.6532e-09

   CompressorIn_bh30_41_81 <= heap_bh30_w19_0 & heap_bh30_w19_7 & heap_bh30_w19_6;
   CompressorIn_bh30_41_82 <= heap_bh30_w20_8 & heap_bh30_w20_7;
      Compressor_bh30_41: Compressor_23_3
      port map ( R => CompressorOut_bh30_41_41,
                 X0 => CompressorIn_bh30_41_81,
                 X1 => CompressorIn_bh30_41_82);
   heap_bh30_w19_8 <= CompressorOut_bh30_41_41(0); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w20_9 <= CompressorOut_bh30_41_41(1); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w21_9 <= CompressorOut_bh30_41_41(2); -- cycle= 0 cp= 1.6532e-09

   CompressorIn_bh30_42_83 <= heap_bh30_w22_0 & heap_bh30_w22_7 & heap_bh30_w22_6;
   CompressorIn_bh30_42_84 <= heap_bh30_w23_9 & heap_bh30_w23_8;
      Compressor_bh30_42: Compressor_23_3
      port map ( R => CompressorOut_bh30_42_42,
                 X0 => CompressorIn_bh30_42_83,
                 X1 => CompressorIn_bh30_42_84);
   heap_bh30_w22_8 <= CompressorOut_bh30_42_42(0); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w23_10 <= CompressorOut_bh30_42_42(1); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w24_10 <= CompressorOut_bh30_42_42(2); -- cycle= 0 cp= 1.6532e-09

   CompressorIn_bh30_43_85 <= heap_bh30_w25_0 & heap_bh30_w25_8 & heap_bh30_w25_7;
   CompressorIn_bh30_43_86 <= heap_bh30_w26_9 & heap_bh30_w26_8;
      Compressor_bh30_43: Compressor_23_3
      port map ( R => CompressorOut_bh30_43_43,
                 X0 => CompressorIn_bh30_43_85,
                 X1 => CompressorIn_bh30_43_86);
   heap_bh30_w25_9 <= CompressorOut_bh30_43_43(0); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w26_10 <= CompressorOut_bh30_43_43(1); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w27_10 <= CompressorOut_bh30_43_43(2); -- cycle= 0 cp= 1.6532e-09

   CompressorIn_bh30_44_87 <= heap_bh30_w28_0 & heap_bh30_w28_8 & heap_bh30_w28_7;
   CompressorIn_bh30_44_88 <= heap_bh30_w29_9 & heap_bh30_w29_8;
      Compressor_bh30_44: Compressor_23_3
      port map ( R => CompressorOut_bh30_44_44,
                 X0 => CompressorIn_bh30_44_87,
                 X1 => CompressorIn_bh30_44_88);
   heap_bh30_w28_9 <= CompressorOut_bh30_44_44(0); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w29_10 <= CompressorOut_bh30_44_44(1); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w30_10 <= CompressorOut_bh30_44_44(2); -- cycle= 0 cp= 1.6532e-09

   CompressorIn_bh30_45_89 <= heap_bh30_w31_0 & heap_bh30_w31_8 & heap_bh30_w31_7;
   CompressorIn_bh30_45_90 <= heap_bh30_w32_9 & heap_bh30_w32_8;
      Compressor_bh30_45: Compressor_23_3
      port map ( R => CompressorOut_bh30_45_45,
                 X0 => CompressorIn_bh30_45_89,
                 X1 => CompressorIn_bh30_45_90);
   heap_bh30_w31_9 <= CompressorOut_bh30_45_45(0); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w32_10 <= CompressorOut_bh30_45_45(1); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w33_10 <= CompressorOut_bh30_45_45(2); -- cycle= 0 cp= 1.6532e-09

   CompressorIn_bh30_46_91 <= heap_bh30_w34_0 & heap_bh30_w34_8 & heap_bh30_w34_7;
   CompressorIn_bh30_46_92 <= heap_bh30_w35_9 & heap_bh30_w35_8;
      Compressor_bh30_46: Compressor_23_3
      port map ( R => CompressorOut_bh30_46_46,
                 X0 => CompressorIn_bh30_46_91,
                 X1 => CompressorIn_bh30_46_92);
   heap_bh30_w34_9 <= CompressorOut_bh30_46_46(0); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w35_10 <= CompressorOut_bh30_46_46(1); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w36_10 <= CompressorOut_bh30_46_46(2); -- cycle= 0 cp= 1.6532e-09

   CompressorIn_bh30_47_93 <= heap_bh30_w37_0 & heap_bh30_w37_9 & heap_bh30_w37_8;
   CompressorIn_bh30_47_94 <= heap_bh30_w38_10 & heap_bh30_w38_9;
      Compressor_bh30_47: Compressor_23_3
      port map ( R => CompressorOut_bh30_47_47,
                 X0 => CompressorIn_bh30_47_93,
                 X1 => CompressorIn_bh30_47_94);
   heap_bh30_w37_10 <= CompressorOut_bh30_47_47(0); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w38_11 <= CompressorOut_bh30_47_47(1); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w39_11 <= CompressorOut_bh30_47_47(2); -- cycle= 0 cp= 1.6532e-09

   CompressorIn_bh30_48_95 <= heap_bh30_w40_0 & heap_bh30_w40_9 & heap_bh30_w40_8;
   CompressorIn_bh30_48_96 <= heap_bh30_w41_10 & heap_bh30_w41_9;
      Compressor_bh30_48: Compressor_23_3
      port map ( R => CompressorOut_bh30_48_48,
                 X0 => CompressorIn_bh30_48_95,
                 X1 => CompressorIn_bh30_48_96);
   heap_bh30_w40_10 <= CompressorOut_bh30_48_48(0); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w41_11 <= CompressorOut_bh30_48_48(1); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w42_11 <= CompressorOut_bh30_48_48(2); -- cycle= 0 cp= 1.6532e-09

   CompressorIn_bh30_49_97 <= heap_bh30_w43_0 & heap_bh30_w43_9 & heap_bh30_w43_8;
   CompressorIn_bh30_49_98 <= heap_bh30_w44_10 & heap_bh30_w44_9;
      Compressor_bh30_49: Compressor_23_3
      port map ( R => CompressorOut_bh30_49_49,
                 X0 => CompressorIn_bh30_49_97,
                 X1 => CompressorIn_bh30_49_98);
   heap_bh30_w43_10 <= CompressorOut_bh30_49_49(0); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w44_11 <= CompressorOut_bh30_49_49(1); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w45_11 <= CompressorOut_bh30_49_49(2); -- cycle= 0 cp= 1.6532e-09

   CompressorIn_bh30_50_99 <= heap_bh30_w46_0 & heap_bh30_w46_9 & heap_bh30_w46_8;
   CompressorIn_bh30_50_100 <= heap_bh30_w47_10 & heap_bh30_w47_9;
      Compressor_bh30_50: Compressor_23_3
      port map ( R => CompressorOut_bh30_50_50,
                 X0 => CompressorIn_bh30_50_99,
                 X1 => CompressorIn_bh30_50_100);
   heap_bh30_w46_10 <= CompressorOut_bh30_50_50(0); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w47_11 <= CompressorOut_bh30_50_50(1); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w48_11 <= CompressorOut_bh30_50_50(2); -- cycle= 0 cp= 1.6532e-09

   CompressorIn_bh30_51_101 <= heap_bh30_w49_0 & heap_bh30_w49_9 & heap_bh30_w49_8;
   CompressorIn_bh30_51_102 <= heap_bh30_w50_10 & heap_bh30_w50_9;
      Compressor_bh30_51: Compressor_23_3
      port map ( R => CompressorOut_bh30_51_51,
                 X0 => CompressorIn_bh30_51_101,
                 X1 => CompressorIn_bh30_51_102);
   heap_bh30_w49_10 <= CompressorOut_bh30_51_51(0); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w50_11 <= CompressorOut_bh30_51_51(1); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w51_11 <= CompressorOut_bh30_51_51(2); -- cycle= 0 cp= 1.6532e-09

   CompressorIn_bh30_52_103 <= heap_bh30_w52_0 & heap_bh30_w52_9 & heap_bh30_w52_8;
   CompressorIn_bh30_52_104 <= heap_bh30_w53_10 & heap_bh30_w53_9;
      Compressor_bh30_52: Compressor_23_3
      port map ( R => CompressorOut_bh30_52_52,
                 X0 => CompressorIn_bh30_52_103,
                 X1 => CompressorIn_bh30_52_104);
   heap_bh30_w52_10 <= CompressorOut_bh30_52_52(0); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w53_11 <= CompressorOut_bh30_52_52(1); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w54_11 <= CompressorOut_bh30_52_52(2); -- cycle= 0 cp= 1.6532e-09

   CompressorIn_bh30_53_105 <= heap_bh30_w55_0 & heap_bh30_w55_9 & heap_bh30_w55_8;
   CompressorIn_bh30_53_106 <= heap_bh30_w56_9 & heap_bh30_w56_8;
      Compressor_bh30_53: Compressor_23_3
      port map ( R => CompressorOut_bh30_53_53,
                 X0 => CompressorIn_bh30_53_105,
                 X1 => CompressorIn_bh30_53_106);
   heap_bh30_w55_10 <= CompressorOut_bh30_53_53(0); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w56_10 <= CompressorOut_bh30_53_53(1); -- cycle= 0 cp= 1.6532e-09
   heap_bh30_w57_9 <= CompressorOut_bh30_53_53(2); -- cycle= 0 cp= 1.6532e-09

   CompressorIn_bh30_54_107 <= heap_bh30_w57_0 & heap_bh30_w57_8 & heap_bh30_w57_9;
   CompressorIn_bh30_54_108 <= heap_bh30_w58_0 & heap_bh30_w58_6;
      Compressor_bh30_54: Compressor_23_3
      port map ( R => CompressorOut_bh30_54_54,
                 X0 => CompressorIn_bh30_54_107,
                 X1 => CompressorIn_bh30_54_108);
   heap_bh30_w57_10 <= CompressorOut_bh30_54_54(0); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w58_7 <= CompressorOut_bh30_54_54(1); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w59_6 <= CompressorOut_bh30_54_54(2); -- cycle= 0 cp= 2.18392e-09

   CompressorIn_bh30_55_109 <= heap_bh30_w9_7 & heap_bh30_w9_6 & heap_bh30_w9_8;
   CompressorIn_bh30_55_110(0) <= heap_bh30_w10_7;
      Compressor_bh30_55: Compressor_13_3
      port map ( R => CompressorOut_bh30_55_55,
                 X0 => CompressorIn_bh30_55_109,
                 X1 => CompressorIn_bh30_55_110);
   heap_bh30_w9_9 <= CompressorOut_bh30_55_55(0); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w10_8 <= CompressorOut_bh30_55_55(1); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w11_9 <= CompressorOut_bh30_55_55(2); -- cycle= 0 cp= 2.18392e-09

   CompressorIn_bh30_56_111 <= heap_bh30_w12_7 & heap_bh30_w12_6 & heap_bh30_w12_8;
   CompressorIn_bh30_56_112(0) <= heap_bh30_w13_8;
      Compressor_bh30_56: Compressor_13_3
      port map ( R => CompressorOut_bh30_56_56,
                 X0 => CompressorIn_bh30_56_111,
                 X1 => CompressorIn_bh30_56_112);
   heap_bh30_w12_9 <= CompressorOut_bh30_56_56(0); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w13_9 <= CompressorOut_bh30_56_56(1); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w14_10 <= CompressorOut_bh30_56_56(2); -- cycle= 0 cp= 2.18392e-09

   CompressorIn_bh30_57_113 <= heap_bh30_w15_8 & heap_bh30_w15_7 & heap_bh30_w15_9;
   CompressorIn_bh30_57_114(0) <= heap_bh30_w16_8;
      Compressor_bh30_57: Compressor_13_3
      port map ( R => CompressorOut_bh30_57_57,
                 X0 => CompressorIn_bh30_57_113,
                 X1 => CompressorIn_bh30_57_114);
   heap_bh30_w15_10 <= CompressorOut_bh30_57_57(0); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w16_9 <= CompressorOut_bh30_57_57(1); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w17_10 <= CompressorOut_bh30_57_57(2); -- cycle= 0 cp= 2.18392e-09

   CompressorIn_bh30_58_115 <= heap_bh30_w18_8 & heap_bh30_w18_7 & heap_bh30_w18_9;
   CompressorIn_bh30_58_116(0) <= heap_bh30_w19_8;
      Compressor_bh30_58: Compressor_13_3
      port map ( R => CompressorOut_bh30_58_58,
                 X0 => CompressorIn_bh30_58_115,
                 X1 => CompressorIn_bh30_58_116);
   heap_bh30_w18_10 <= CompressorOut_bh30_58_58(0); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w19_9 <= CompressorOut_bh30_58_58(1); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w20_10 <= CompressorOut_bh30_58_58(2); -- cycle= 0 cp= 2.18392e-09

   CompressorIn_bh30_59_117 <= heap_bh30_w21_8 & heap_bh30_w21_7 & heap_bh30_w21_9;
   CompressorIn_bh30_59_118(0) <= heap_bh30_w22_8;
      Compressor_bh30_59: Compressor_13_3
      port map ( R => CompressorOut_bh30_59_59,
                 X0 => CompressorIn_bh30_59_117,
                 X1 => CompressorIn_bh30_59_118);
   heap_bh30_w21_10 <= CompressorOut_bh30_59_59(0); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w22_9 <= CompressorOut_bh30_59_59(1); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w23_11 <= CompressorOut_bh30_59_59(2); -- cycle= 0 cp= 2.18392e-09

   CompressorIn_bh30_60_119 <= heap_bh30_w24_9 & heap_bh30_w24_8 & heap_bh30_w24_10;
   CompressorIn_bh30_60_120(0) <= heap_bh30_w25_9;
      Compressor_bh30_60: Compressor_13_3
      port map ( R => CompressorOut_bh30_60_60,
                 X0 => CompressorIn_bh30_60_119,
                 X1 => CompressorIn_bh30_60_120);
   heap_bh30_w24_11 <= CompressorOut_bh30_60_60(0); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w25_10 <= CompressorOut_bh30_60_60(1); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w26_11 <= CompressorOut_bh30_60_60(2); -- cycle= 0 cp= 2.18392e-09

   CompressorIn_bh30_61_121 <= heap_bh30_w27_9 & heap_bh30_w27_8 & heap_bh30_w27_10;
   CompressorIn_bh30_61_122(0) <= heap_bh30_w28_9;
      Compressor_bh30_61: Compressor_13_3
      port map ( R => CompressorOut_bh30_61_61,
                 X0 => CompressorIn_bh30_61_121,
                 X1 => CompressorIn_bh30_61_122);
   heap_bh30_w27_11 <= CompressorOut_bh30_61_61(0); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w28_10 <= CompressorOut_bh30_61_61(1); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w29_11 <= CompressorOut_bh30_61_61(2); -- cycle= 0 cp= 2.18392e-09

   CompressorIn_bh30_62_123 <= heap_bh30_w30_9 & heap_bh30_w30_8 & heap_bh30_w30_10;
   CompressorIn_bh30_62_124(0) <= heap_bh30_w31_9;
      Compressor_bh30_62: Compressor_13_3
      port map ( R => CompressorOut_bh30_62_62,
                 X0 => CompressorIn_bh30_62_123,
                 X1 => CompressorIn_bh30_62_124);
   heap_bh30_w30_11 <= CompressorOut_bh30_62_62(0); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w31_10 <= CompressorOut_bh30_62_62(1); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w32_11 <= CompressorOut_bh30_62_62(2); -- cycle= 0 cp= 2.18392e-09

   CompressorIn_bh30_63_125 <= heap_bh30_w33_9 & heap_bh30_w33_8 & heap_bh30_w33_10;
   CompressorIn_bh30_63_126(0) <= heap_bh30_w34_9;
      Compressor_bh30_63: Compressor_13_3
      port map ( R => CompressorOut_bh30_63_63,
                 X0 => CompressorIn_bh30_63_125,
                 X1 => CompressorIn_bh30_63_126);
   heap_bh30_w33_11 <= CompressorOut_bh30_63_63(0); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w34_10 <= CompressorOut_bh30_63_63(1); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w35_11 <= CompressorOut_bh30_63_63(2); -- cycle= 0 cp= 2.18392e-09

   CompressorIn_bh30_64_127 <= heap_bh30_w36_9 & heap_bh30_w36_8 & heap_bh30_w36_10;
   CompressorIn_bh30_64_128(0) <= heap_bh30_w37_10;
      Compressor_bh30_64: Compressor_13_3
      port map ( R => CompressorOut_bh30_64_64,
                 X0 => CompressorIn_bh30_64_127,
                 X1 => CompressorIn_bh30_64_128);
   heap_bh30_w36_11 <= CompressorOut_bh30_64_64(0); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w37_11 <= CompressorOut_bh30_64_64(1); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w38_12 <= CompressorOut_bh30_64_64(2); -- cycle= 0 cp= 2.18392e-09

   CompressorIn_bh30_65_129 <= heap_bh30_w39_10 & heap_bh30_w39_9 & heap_bh30_w39_11;
   CompressorIn_bh30_65_130(0) <= heap_bh30_w40_10;
      Compressor_bh30_65: Compressor_13_3
      port map ( R => CompressorOut_bh30_65_65,
                 X0 => CompressorIn_bh30_65_129,
                 X1 => CompressorIn_bh30_65_130);
   heap_bh30_w39_12 <= CompressorOut_bh30_65_65(0); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w40_11 <= CompressorOut_bh30_65_65(1); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w41_12 <= CompressorOut_bh30_65_65(2); -- cycle= 0 cp= 2.18392e-09

   CompressorIn_bh30_66_131 <= heap_bh30_w42_10 & heap_bh30_w42_9 & heap_bh30_w42_11;
   CompressorIn_bh30_66_132(0) <= heap_bh30_w43_10;
      Compressor_bh30_66: Compressor_13_3
      port map ( R => CompressorOut_bh30_66_66,
                 X0 => CompressorIn_bh30_66_131,
                 X1 => CompressorIn_bh30_66_132);
   heap_bh30_w42_12 <= CompressorOut_bh30_66_66(0); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w43_11 <= CompressorOut_bh30_66_66(1); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w44_12 <= CompressorOut_bh30_66_66(2); -- cycle= 0 cp= 2.18392e-09

   CompressorIn_bh30_67_133 <= heap_bh30_w45_10 & heap_bh30_w45_9 & heap_bh30_w45_11;
   CompressorIn_bh30_67_134(0) <= heap_bh30_w46_10;
      Compressor_bh30_67: Compressor_13_3
      port map ( R => CompressorOut_bh30_67_67,
                 X0 => CompressorIn_bh30_67_133,
                 X1 => CompressorIn_bh30_67_134);
   heap_bh30_w45_12 <= CompressorOut_bh30_67_67(0); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w46_11 <= CompressorOut_bh30_67_67(1); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w47_12 <= CompressorOut_bh30_67_67(2); -- cycle= 0 cp= 2.18392e-09

   CompressorIn_bh30_68_135 <= heap_bh30_w48_10 & heap_bh30_w48_9 & heap_bh30_w48_11;
   CompressorIn_bh30_68_136(0) <= heap_bh30_w49_10;
      Compressor_bh30_68: Compressor_13_3
      port map ( R => CompressorOut_bh30_68_68,
                 X0 => CompressorIn_bh30_68_135,
                 X1 => CompressorIn_bh30_68_136);
   heap_bh30_w48_12 <= CompressorOut_bh30_68_68(0); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w49_11 <= CompressorOut_bh30_68_68(1); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w50_12 <= CompressorOut_bh30_68_68(2); -- cycle= 0 cp= 2.18392e-09

   CompressorIn_bh30_69_137 <= heap_bh30_w51_10 & heap_bh30_w51_9 & heap_bh30_w51_11;
   CompressorIn_bh30_69_138(0) <= heap_bh30_w52_10;
      Compressor_bh30_69: Compressor_13_3
      port map ( R => CompressorOut_bh30_69_69,
                 X0 => CompressorIn_bh30_69_137,
                 X1 => CompressorIn_bh30_69_138);
   heap_bh30_w51_12 <= CompressorOut_bh30_69_69(0); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w52_11 <= CompressorOut_bh30_69_69(1); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w53_12 <= CompressorOut_bh30_69_69(2); -- cycle= 0 cp= 2.18392e-09

   CompressorIn_bh30_70_139 <= heap_bh30_w54_10 & heap_bh30_w54_9 & heap_bh30_w54_11;
   CompressorIn_bh30_70_140(0) <= heap_bh30_w55_10;
      Compressor_bh30_70: Compressor_13_3
      port map ( R => CompressorOut_bh30_70_70,
                 X0 => CompressorIn_bh30_70_139,
                 X1 => CompressorIn_bh30_70_140);
   heap_bh30_w54_12 <= CompressorOut_bh30_70_70(0); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w55_11 <= CompressorOut_bh30_70_70(1); -- cycle= 0 cp= 2.18392e-09
   heap_bh30_w56_11 <= CompressorOut_bh30_70_70(2); -- cycle= 0 cp= 2.18392e-09

   CompressorIn_bh30_71_141 <= heap_bh30_w23_10 & heap_bh30_w23_11 & heap_bh30_w23_7 & heap_bh30_w23_6 & heap_bh30_w23_5 & heap_bh30_w23_4;
      Compressor_bh30_71: Compressor_6_3
      port map ( R => CompressorOut_bh30_71_71,
                 X0 => CompressorIn_bh30_71_141);
   heap_bh30_w23_12 <= CompressorOut_bh30_71_71(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w24_12 <= CompressorOut_bh30_71_71(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w25_11 <= CompressorOut_bh30_71_71(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_72_142 <= heap_bh30_w26_10 & heap_bh30_w26_11 & heap_bh30_w26_7 & heap_bh30_w26_6 & heap_bh30_w26_5 & heap_bh30_w26_4;
      Compressor_bh30_72: Compressor_6_3
      port map ( R => CompressorOut_bh30_72_72,
                 X0 => CompressorIn_bh30_72_142);
   heap_bh30_w26_12 <= CompressorOut_bh30_72_72(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w27_12 <= CompressorOut_bh30_72_72(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w28_11 <= CompressorOut_bh30_72_72(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_73_143 <= heap_bh30_w29_10 & heap_bh30_w29_11 & heap_bh30_w29_7 & heap_bh30_w29_6 & heap_bh30_w29_5 & heap_bh30_w29_4;
      Compressor_bh30_73: Compressor_6_3
      port map ( R => CompressorOut_bh30_73_73,
                 X0 => CompressorIn_bh30_73_143);
   heap_bh30_w29_12 <= CompressorOut_bh30_73_73(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w30_12 <= CompressorOut_bh30_73_73(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w31_11 <= CompressorOut_bh30_73_73(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_74_144 <= heap_bh30_w32_10 & heap_bh30_w32_11 & heap_bh30_w32_7 & heap_bh30_w32_6 & heap_bh30_w32_5 & heap_bh30_w32_4;
      Compressor_bh30_74: Compressor_6_3
      port map ( R => CompressorOut_bh30_74_74,
                 X0 => CompressorIn_bh30_74_144);
   heap_bh30_w32_12 <= CompressorOut_bh30_74_74(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w33_12 <= CompressorOut_bh30_74_74(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w34_11 <= CompressorOut_bh30_74_74(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_75_145 <= heap_bh30_w35_10 & heap_bh30_w35_11 & heap_bh30_w35_7 & heap_bh30_w35_6 & heap_bh30_w35_5 & heap_bh30_w35_4;
      Compressor_bh30_75: Compressor_6_3
      port map ( R => CompressorOut_bh30_75_75,
                 X0 => CompressorIn_bh30_75_145);
   heap_bh30_w35_12 <= CompressorOut_bh30_75_75(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w36_12 <= CompressorOut_bh30_75_75(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w37_12 <= CompressorOut_bh30_75_75(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_76_146 <= heap_bh30_w37_11 & heap_bh30_w37_7 & heap_bh30_w37_6 & heap_bh30_w37_5 & heap_bh30_w37_4 & heap_bh30_w37_3;
      Compressor_bh30_76: Compressor_6_3
      port map ( R => CompressorOut_bh30_76_76,
                 X0 => CompressorIn_bh30_76_146);
   heap_bh30_w37_13 <= CompressorOut_bh30_76_76(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w38_13 <= CompressorOut_bh30_76_76(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w39_13 <= CompressorOut_bh30_76_76(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_77_147 <= heap_bh30_w38_11 & heap_bh30_w38_12 & heap_bh30_w38_8 & heap_bh30_w38_7 & heap_bh30_w38_6 & heap_bh30_w38_5;
      Compressor_bh30_77: Compressor_6_3
      port map ( R => CompressorOut_bh30_77_77,
                 X0 => CompressorIn_bh30_77_147);
   heap_bh30_w38_14 <= CompressorOut_bh30_77_77(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w39_14 <= CompressorOut_bh30_77_77(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w40_12 <= CompressorOut_bh30_77_77(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_78_148 <= heap_bh30_w39_12 & heap_bh30_w39_8 & heap_bh30_w39_7 & heap_bh30_w39_6 & heap_bh30_w39_5 & heap_bh30_w39_4;
      Compressor_bh30_78: Compressor_6_3
      port map ( R => CompressorOut_bh30_78_78,
                 X0 => CompressorIn_bh30_78_148);
   heap_bh30_w39_15 <= CompressorOut_bh30_78_78(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w40_13 <= CompressorOut_bh30_78_78(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w41_13 <= CompressorOut_bh30_78_78(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_79_149 <= heap_bh30_w40_11 & heap_bh30_w40_7 & heap_bh30_w40_6 & heap_bh30_w40_5 & heap_bh30_w40_4 & heap_bh30_w40_3;
      Compressor_bh30_79: Compressor_6_3
      port map ( R => CompressorOut_bh30_79_79,
                 X0 => CompressorIn_bh30_79_149);
   heap_bh30_w40_14 <= CompressorOut_bh30_79_79(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w41_14 <= CompressorOut_bh30_79_79(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w42_13 <= CompressorOut_bh30_79_79(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_80_150 <= heap_bh30_w41_11 & heap_bh30_w41_12 & heap_bh30_w41_8 & heap_bh30_w41_7 & heap_bh30_w41_6 & heap_bh30_w41_5;
      Compressor_bh30_80: Compressor_6_3
      port map ( R => CompressorOut_bh30_80_80,
                 X0 => CompressorIn_bh30_80_150);
   heap_bh30_w41_15 <= CompressorOut_bh30_80_80(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w42_14 <= CompressorOut_bh30_80_80(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w43_12 <= CompressorOut_bh30_80_80(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_81_151 <= heap_bh30_w42_12 & heap_bh30_w42_8 & heap_bh30_w42_7 & heap_bh30_w42_6 & heap_bh30_w42_5 & heap_bh30_w42_4;
      Compressor_bh30_81: Compressor_6_3
      port map ( R => CompressorOut_bh30_81_81,
                 X0 => CompressorIn_bh30_81_151);
   heap_bh30_w42_15 <= CompressorOut_bh30_81_81(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w43_13 <= CompressorOut_bh30_81_81(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w44_13 <= CompressorOut_bh30_81_81(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_82_152 <= heap_bh30_w43_11 & heap_bh30_w43_7 & heap_bh30_w43_6 & heap_bh30_w43_5 & heap_bh30_w43_4 & heap_bh30_w43_3;
      Compressor_bh30_82: Compressor_6_3
      port map ( R => CompressorOut_bh30_82_82,
                 X0 => CompressorIn_bh30_82_152);
   heap_bh30_w43_14 <= CompressorOut_bh30_82_82(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w44_14 <= CompressorOut_bh30_82_82(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w45_13 <= CompressorOut_bh30_82_82(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_83_153 <= heap_bh30_w44_11 & heap_bh30_w44_12 & heap_bh30_w44_8 & heap_bh30_w44_7 & heap_bh30_w44_6 & heap_bh30_w44_5;
      Compressor_bh30_83: Compressor_6_3
      port map ( R => CompressorOut_bh30_83_83,
                 X0 => CompressorIn_bh30_83_153);
   heap_bh30_w44_15 <= CompressorOut_bh30_83_83(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w45_14 <= CompressorOut_bh30_83_83(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w46_12 <= CompressorOut_bh30_83_83(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_84_154 <= heap_bh30_w45_12 & heap_bh30_w45_8 & heap_bh30_w45_7 & heap_bh30_w45_6 & heap_bh30_w45_5 & heap_bh30_w45_4;
      Compressor_bh30_84: Compressor_6_3
      port map ( R => CompressorOut_bh30_84_84,
                 X0 => CompressorIn_bh30_84_154);
   heap_bh30_w45_15 <= CompressorOut_bh30_84_84(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w46_13 <= CompressorOut_bh30_84_84(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w47_13 <= CompressorOut_bh30_84_84(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_85_155 <= heap_bh30_w46_11 & heap_bh30_w46_7 & heap_bh30_w46_6 & heap_bh30_w46_5 & heap_bh30_w46_4 & heap_bh30_w46_3;
      Compressor_bh30_85: Compressor_6_3
      port map ( R => CompressorOut_bh30_85_85,
                 X0 => CompressorIn_bh30_85_155);
   heap_bh30_w46_14 <= CompressorOut_bh30_85_85(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w47_14 <= CompressorOut_bh30_85_85(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w48_13 <= CompressorOut_bh30_85_85(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_86_156 <= heap_bh30_w47_11 & heap_bh30_w47_12 & heap_bh30_w47_8 & heap_bh30_w47_7 & heap_bh30_w47_6 & heap_bh30_w47_5;
      Compressor_bh30_86: Compressor_6_3
      port map ( R => CompressorOut_bh30_86_86,
                 X0 => CompressorIn_bh30_86_156);
   heap_bh30_w47_15 <= CompressorOut_bh30_86_86(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w48_14 <= CompressorOut_bh30_86_86(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w49_12 <= CompressorOut_bh30_86_86(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_87_157 <= heap_bh30_w48_12 & heap_bh30_w48_8 & heap_bh30_w48_7 & heap_bh30_w48_6 & heap_bh30_w48_5 & heap_bh30_w48_4;
      Compressor_bh30_87: Compressor_6_3
      port map ( R => CompressorOut_bh30_87_87,
                 X0 => CompressorIn_bh30_87_157);
   heap_bh30_w48_15 <= CompressorOut_bh30_87_87(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w49_13 <= CompressorOut_bh30_87_87(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w50_13 <= CompressorOut_bh30_87_87(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_88_158 <= heap_bh30_w49_11 & heap_bh30_w49_7 & heap_bh30_w49_6 & heap_bh30_w49_5 & heap_bh30_w49_4 & heap_bh30_w49_3;
      Compressor_bh30_88: Compressor_6_3
      port map ( R => CompressorOut_bh30_88_88,
                 X0 => CompressorIn_bh30_88_158);
   heap_bh30_w49_14 <= CompressorOut_bh30_88_88(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w50_14 <= CompressorOut_bh30_88_88(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w51_13 <= CompressorOut_bh30_88_88(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_89_159 <= heap_bh30_w50_11 & heap_bh30_w50_12 & heap_bh30_w50_8 & heap_bh30_w50_7 & heap_bh30_w50_6 & heap_bh30_w50_5;
      Compressor_bh30_89: Compressor_6_3
      port map ( R => CompressorOut_bh30_89_89,
                 X0 => CompressorIn_bh30_89_159);
   heap_bh30_w50_15 <= CompressorOut_bh30_89_89(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w51_14 <= CompressorOut_bh30_89_89(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w52_12 <= CompressorOut_bh30_89_89(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_90_160 <= heap_bh30_w51_12 & heap_bh30_w51_8 & heap_bh30_w51_7 & heap_bh30_w51_6 & heap_bh30_w51_5 & heap_bh30_w51_4;
      Compressor_bh30_90: Compressor_6_3
      port map ( R => CompressorOut_bh30_90_90,
                 X0 => CompressorIn_bh30_90_160);
   heap_bh30_w51_15 <= CompressorOut_bh30_90_90(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w52_13 <= CompressorOut_bh30_90_90(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w53_13 <= CompressorOut_bh30_90_90(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_91_161 <= heap_bh30_w52_11 & heap_bh30_w52_7 & heap_bh30_w52_6 & heap_bh30_w52_5 & heap_bh30_w52_4 & heap_bh30_w52_3;
      Compressor_bh30_91: Compressor_6_3
      port map ( R => CompressorOut_bh30_91_91,
                 X0 => CompressorIn_bh30_91_161);
   heap_bh30_w52_14 <= CompressorOut_bh30_91_91(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w53_14 <= CompressorOut_bh30_91_91(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w54_13 <= CompressorOut_bh30_91_91(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_92_162 <= heap_bh30_w53_11 & heap_bh30_w53_12 & heap_bh30_w53_8 & heap_bh30_w53_7 & heap_bh30_w53_6 & heap_bh30_w53_5;
      Compressor_bh30_92: Compressor_6_3
      port map ( R => CompressorOut_bh30_92_92,
                 X0 => CompressorIn_bh30_92_162);
   heap_bh30_w53_15 <= CompressorOut_bh30_92_92(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w54_14 <= CompressorOut_bh30_92_92(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w55_12 <= CompressorOut_bh30_92_92(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_93_163 <= heap_bh30_w54_12 & heap_bh30_w54_8 & heap_bh30_w54_7 & heap_bh30_w54_6 & heap_bh30_w54_5 & heap_bh30_w54_4;
      Compressor_bh30_93: Compressor_6_3
      port map ( R => CompressorOut_bh30_93_93,
                 X0 => CompressorIn_bh30_93_163);
   heap_bh30_w54_15 <= CompressorOut_bh30_93_93(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w55_13 <= CompressorOut_bh30_93_93(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w56_12 <= CompressorOut_bh30_93_93(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_94_164 <= heap_bh30_w55_11 & heap_bh30_w55_7 & heap_bh30_w55_6 & heap_bh30_w55_5 & heap_bh30_w55_4 & heap_bh30_w55_3;
      Compressor_bh30_94: Compressor_6_3
      port map ( R => CompressorOut_bh30_94_94,
                 X0 => CompressorIn_bh30_94_164);
   heap_bh30_w55_14 <= CompressorOut_bh30_94_94(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w56_13 <= CompressorOut_bh30_94_94(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w57_11 <= CompressorOut_bh30_94_94(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_95_165 <= heap_bh30_w56_10 & heap_bh30_w56_11 & heap_bh30_w56_7 & heap_bh30_w56_6 & heap_bh30_w56_5 & heap_bh30_w56_4;
      Compressor_bh30_95: Compressor_6_3
      port map ( R => CompressorOut_bh30_95_95,
                 X0 => CompressorIn_bh30_95_165);
   heap_bh30_w56_14 <= CompressorOut_bh30_95_95(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w57_12 <= CompressorOut_bh30_95_95(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w58_8 <= CompressorOut_bh30_95_95(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_96_166 <= heap_bh30_w57_10 & heap_bh30_w57_7 & heap_bh30_w57_6 & heap_bh30_w57_5 & heap_bh30_w57_4 & heap_bh30_w57_3;
      Compressor_bh30_96: Compressor_6_3
      port map ( R => CompressorOut_bh30_96_96,
                 X0 => CompressorIn_bh30_96_166);
   heap_bh30_w57_13 <= CompressorOut_bh30_96_96(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w58_9 <= CompressorOut_bh30_96_96(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w59_7 <= CompressorOut_bh30_96_96(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_97_167 <= heap_bh30_w58_7 & heap_bh30_w58_5 & heap_bh30_w58_4 & heap_bh30_w58_3 & heap_bh30_w58_2 & heap_bh30_w58_1;
      Compressor_bh30_97: Compressor_6_3
      port map ( R => CompressorOut_bh30_97_97,
                 X0 => CompressorIn_bh30_97_167);
   heap_bh30_w58_10 <= CompressorOut_bh30_97_97(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w59_8 <= CompressorOut_bh30_97_97(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w60_6 <= CompressorOut_bh30_97_97(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_98_168 <= heap_bh30_w59_0 & heap_bh30_w59_6 & heap_bh30_w59_5 & heap_bh30_w59_4 & heap_bh30_w59_3 & heap_bh30_w59_2;
      Compressor_bh30_98: Compressor_6_3
      port map ( R => CompressorOut_bh30_98_98,
                 X0 => CompressorIn_bh30_98_168);
   heap_bh30_w59_9 <= CompressorOut_bh30_98_98(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w60_7 <= CompressorOut_bh30_98_98(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w61_5 <= CompressorOut_bh30_98_98(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_99_169 <= heap_bh30_w60_0 & heap_bh30_w60_5 & heap_bh30_w60_4 & heap_bh30_w60_3 & heap_bh30_w60_2 & heap_bh30_w60_1;
      Compressor_bh30_99: Compressor_6_3
      port map ( R => CompressorOut_bh30_99_99,
                 X0 => CompressorIn_bh30_99_169);
   heap_bh30_w60_8 <= CompressorOut_bh30_99_99(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w61_6 <= CompressorOut_bh30_99_99(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w62_5 <= CompressorOut_bh30_99_99(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_100_170 <= heap_bh30_w6_7 & heap_bh30_w6_6 & heap_bh30_w6_5 & heap_bh30_w6_4;
   CompressorIn_bh30_100_171(0) <= heap_bh30_w7_7;
      Compressor_bh30_100: Compressor_14_3
      port map ( R => CompressorOut_bh30_100_100,
                 X0 => CompressorIn_bh30_100_170,
                 X1 => CompressorIn_bh30_100_171);
   heap_bh30_w6_8 <= CompressorOut_bh30_100_100(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w7_8 <= CompressorOut_bh30_100_100(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w8_9 <= CompressorOut_bh30_100_100(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_101_172 <= heap_bh30_w11_8 & heap_bh30_w11_9 & heap_bh30_w11_5 & heap_bh30_w11_4;
   CompressorIn_bh30_101_173(0) <= heap_bh30_w12_9;
      Compressor_bh30_101: Compressor_14_3
      port map ( R => CompressorOut_bh30_101_101,
                 X0 => CompressorIn_bh30_101_172,
                 X1 => CompressorIn_bh30_101_173);
   heap_bh30_w11_10 <= CompressorOut_bh30_101_101(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w12_10 <= CompressorOut_bh30_101_101(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w13_10 <= CompressorOut_bh30_101_101(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_102_174 <= heap_bh30_w13_9 & heap_bh30_w13_5 & heap_bh30_w13_4 & heap_bh30_w13_3;
   CompressorIn_bh30_102_175(0) <= heap_bh30_w14_9;
      Compressor_bh30_102: Compressor_14_3
      port map ( R => CompressorOut_bh30_102_102,
                 X0 => CompressorIn_bh30_102_174,
                 X1 => CompressorIn_bh30_102_175);
   heap_bh30_w13_11 <= CompressorOut_bh30_102_102(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w14_11 <= CompressorOut_bh30_102_102(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w15_11 <= CompressorOut_bh30_102_102(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_103_176 <= heap_bh30_w14_10 & heap_bh30_w14_6 & heap_bh30_w14_5 & heap_bh30_w14_4;
   CompressorIn_bh30_103_177(0) <= heap_bh30_w15_10;
      Compressor_bh30_103: Compressor_14_3
      port map ( R => CompressorOut_bh30_103_103,
                 X0 => CompressorIn_bh30_103_176,
                 X1 => CompressorIn_bh30_103_177);
   heap_bh30_w14_12 <= CompressorOut_bh30_103_103(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w15_12 <= CompressorOut_bh30_103_103(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w16_10 <= CompressorOut_bh30_103_103(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_104_178 <= heap_bh30_w16_9 & heap_bh30_w16_5 & heap_bh30_w16_4 & heap_bh30_w16_3;
   CompressorIn_bh30_104_179(0) <= heap_bh30_w17_9;
      Compressor_bh30_104: Compressor_14_3
      port map ( R => CompressorOut_bh30_104_104,
                 X0 => CompressorIn_bh30_104_178,
                 X1 => CompressorIn_bh30_104_179);
   heap_bh30_w16_11 <= CompressorOut_bh30_104_104(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w17_11 <= CompressorOut_bh30_104_104(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w18_11 <= CompressorOut_bh30_104_104(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_105_180 <= heap_bh30_w17_10 & heap_bh30_w17_6 & heap_bh30_w17_5 & heap_bh30_w17_4;
   CompressorIn_bh30_105_181(0) <= heap_bh30_w18_10;
      Compressor_bh30_105: Compressor_14_3
      port map ( R => CompressorOut_bh30_105_105,
                 X0 => CompressorIn_bh30_105_180,
                 X1 => CompressorIn_bh30_105_181);
   heap_bh30_w17_12 <= CompressorOut_bh30_105_105(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w18_12 <= CompressorOut_bh30_105_105(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w19_10 <= CompressorOut_bh30_105_105(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_106_182 <= heap_bh30_w19_9 & heap_bh30_w19_5 & heap_bh30_w19_4 & heap_bh30_w19_3;
   CompressorIn_bh30_106_183(0) <= heap_bh30_w20_9;
      Compressor_bh30_106: Compressor_14_3
      port map ( R => CompressorOut_bh30_106_106,
                 X0 => CompressorIn_bh30_106_182,
                 X1 => CompressorIn_bh30_106_183);
   heap_bh30_w19_11 <= CompressorOut_bh30_106_106(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w20_11 <= CompressorOut_bh30_106_106(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w21_11 <= CompressorOut_bh30_106_106(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_107_184 <= heap_bh30_w20_10 & heap_bh30_w20_6 & heap_bh30_w20_5 & heap_bh30_w20_4;
   CompressorIn_bh30_107_185(0) <= heap_bh30_w21_10;
      Compressor_bh30_107: Compressor_14_3
      port map ( R => CompressorOut_bh30_107_107,
                 X0 => CompressorIn_bh30_107_184,
                 X1 => CompressorIn_bh30_107_185);
   heap_bh30_w20_12 <= CompressorOut_bh30_107_107(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w21_12 <= CompressorOut_bh30_107_107(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w22_10 <= CompressorOut_bh30_107_107(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_108_186 <= heap_bh30_w24_11 & heap_bh30_w24_7 & heap_bh30_w24_6 & heap_bh30_w24_5;
   CompressorIn_bh30_108_187(0) <= heap_bh30_w25_10;
      Compressor_bh30_108: Compressor_14_3
      port map ( R => CompressorOut_bh30_108_108,
                 X0 => CompressorIn_bh30_108_186,
                 X1 => CompressorIn_bh30_108_187);
   heap_bh30_w24_13 <= CompressorOut_bh30_108_108(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w25_12 <= CompressorOut_bh30_108_108(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w26_13 <= CompressorOut_bh30_108_108(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_109_188 <= heap_bh30_w27_11 & heap_bh30_w27_7 & heap_bh30_w27_6 & heap_bh30_w27_5;
   CompressorIn_bh30_109_189(0) <= heap_bh30_w28_10;
      Compressor_bh30_109: Compressor_14_3
      port map ( R => CompressorOut_bh30_109_109,
                 X0 => CompressorIn_bh30_109_188,
                 X1 => CompressorIn_bh30_109_189);
   heap_bh30_w27_13 <= CompressorOut_bh30_109_109(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w28_12 <= CompressorOut_bh30_109_109(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w29_13 <= CompressorOut_bh30_109_109(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_110_190 <= heap_bh30_w30_11 & heap_bh30_w30_7 & heap_bh30_w30_6 & heap_bh30_w30_5;
   CompressorIn_bh30_110_191(0) <= heap_bh30_w31_10;
      Compressor_bh30_110: Compressor_14_3
      port map ( R => CompressorOut_bh30_110_110,
                 X0 => CompressorIn_bh30_110_190,
                 X1 => CompressorIn_bh30_110_191);
   heap_bh30_w30_13 <= CompressorOut_bh30_110_110(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w31_12 <= CompressorOut_bh30_110_110(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w32_13 <= CompressorOut_bh30_110_110(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_111_192 <= heap_bh30_w33_11 & heap_bh30_w33_7 & heap_bh30_w33_6 & heap_bh30_w33_5;
   CompressorIn_bh30_111_193(0) <= heap_bh30_w34_10;
      Compressor_bh30_111: Compressor_14_3
      port map ( R => CompressorOut_bh30_111_111,
                 X0 => CompressorIn_bh30_111_192,
                 X1 => CompressorIn_bh30_111_193);
   heap_bh30_w33_13 <= CompressorOut_bh30_111_111(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w34_12 <= CompressorOut_bh30_111_111(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w35_13 <= CompressorOut_bh30_111_111(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_112_194 <= heap_bh30_w61_4 & heap_bh30_w61_3 & heap_bh30_w61_2 & heap_bh30_w61_1;
   CompressorIn_bh30_112_195(0) <= heap_bh30_w62_4;
      Compressor_bh30_112: Compressor_14_3
      port map ( R => CompressorOut_bh30_112_112,
                 X0 => CompressorIn_bh30_112_194,
                 X1 => CompressorIn_bh30_112_195);
   heap_bh30_w61_7 <= CompressorOut_bh30_112_112(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w62_6 <= CompressorOut_bh30_112_112(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w63_5 <= CompressorOut_bh30_112_112(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_113_196 <= heap_bh30_w62_3 & heap_bh30_w62_2 & heap_bh30_w62_1 & heap_bh30_w62_0;
   CompressorIn_bh30_113_197(0) <= heap_bh30_w63_4;
      Compressor_bh30_113: Compressor_14_3
      port map ( R => CompressorOut_bh30_113_113,
                 X0 => CompressorIn_bh30_113_196,
                 X1 => CompressorIn_bh30_113_197);
   heap_bh30_w62_7 <= CompressorOut_bh30_113_113(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w63_6 <= CompressorOut_bh30_113_113(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w64_4 <= CompressorOut_bh30_113_113(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_114_198 <= heap_bh30_w63_3 & heap_bh30_w63_2 & heap_bh30_w63_1 & heap_bh30_w63_0;
   CompressorIn_bh30_114_199(0) <= heap_bh30_w64_3;
      Compressor_bh30_114: Compressor_14_3
      port map ( R => CompressorOut_bh30_114_114,
                 X0 => CompressorIn_bh30_114_198,
                 X1 => CompressorIn_bh30_114_199);
   heap_bh30_w63_7 <= CompressorOut_bh30_114_114(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w64_5 <= CompressorOut_bh30_114_114(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w65_4 <= CompressorOut_bh30_114_114(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_115_200 <= heap_bh30_w65_3 & heap_bh30_w65_2 & heap_bh30_w65_1 & heap_bh30_w65_0;
   CompressorIn_bh30_115_201(0) <= heap_bh30_w66_3;
      Compressor_bh30_115: Compressor_14_3
      port map ( R => CompressorOut_bh30_115_115,
                 X0 => CompressorIn_bh30_115_200,
                 X1 => CompressorIn_bh30_115_201);
   heap_bh30_w65_5 <= CompressorOut_bh30_115_115(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w66_4 <= CompressorOut_bh30_115_115(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w67_4 <= CompressorOut_bh30_115_115(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_116_202 <= heap_bh30_w67_3 & heap_bh30_w67_2 & heap_bh30_w67_1 & heap_bh30_w67_0;
   CompressorIn_bh30_116_203(0) <= heap_bh30_w68_3;
      Compressor_bh30_116: Compressor_14_3
      port map ( R => CompressorOut_bh30_116_116,
                 X0 => CompressorIn_bh30_116_202,
                 X1 => CompressorIn_bh30_116_203);
   heap_bh30_w67_5 <= CompressorOut_bh30_116_116(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w68_4 <= CompressorOut_bh30_116_116(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w69_4 <= CompressorOut_bh30_116_116(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_117_204 <= heap_bh30_w69_3 & heap_bh30_w69_2 & heap_bh30_w69_1 & heap_bh30_w69_0;
   CompressorIn_bh30_117_205(0) <= heap_bh30_w70_3;
      Compressor_bh30_117: Compressor_14_3
      port map ( R => CompressorOut_bh30_117_117,
                 X0 => CompressorIn_bh30_117_204,
                 X1 => CompressorIn_bh30_117_205);
   heap_bh30_w69_5 <= CompressorOut_bh30_117_117(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w70_4 <= CompressorOut_bh30_117_117(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w71_4 <= CompressorOut_bh30_117_117(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_118_206 <= heap_bh30_w71_3 & heap_bh30_w71_2 & heap_bh30_w71_1 & heap_bh30_w71_0;
   CompressorIn_bh30_118_207(0) <= heap_bh30_w72_3;
      Compressor_bh30_118: Compressor_14_3
      port map ( R => CompressorOut_bh30_118_118,
                 X0 => CompressorIn_bh30_118_206,
                 X1 => CompressorIn_bh30_118_207);
   heap_bh30_w71_5 <= CompressorOut_bh30_118_118(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w72_4 <= CompressorOut_bh30_118_118(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w73_4 <= CompressorOut_bh30_118_118(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_119_208 <= heap_bh30_w73_3 & heap_bh30_w73_2 & heap_bh30_w73_1 & heap_bh30_w73_0;
   CompressorIn_bh30_119_209(0) <= heap_bh30_w74_3;
      Compressor_bh30_119: Compressor_14_3
      port map ( R => CompressorOut_bh30_119_119,
                 X0 => CompressorIn_bh30_119_208,
                 X1 => CompressorIn_bh30_119_209);
   heap_bh30_w73_5 <= CompressorOut_bh30_119_119(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w74_4 <= CompressorOut_bh30_119_119(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w75_4 <= CompressorOut_bh30_119_119(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_120_210 <= heap_bh30_w75_3 & heap_bh30_w75_2 & heap_bh30_w75_1 & heap_bh30_w75_0;
   CompressorIn_bh30_120_211(0) <= heap_bh30_w76_3;
      Compressor_bh30_120: Compressor_14_3
      port map ( R => CompressorOut_bh30_120_120,
                 X0 => CompressorIn_bh30_120_210,
                 X1 => CompressorIn_bh30_120_211);
   heap_bh30_w75_5 <= CompressorOut_bh30_120_120(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w76_4 <= CompressorOut_bh30_120_120(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w77_4 <= CompressorOut_bh30_120_120(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_121_212 <= heap_bh30_w77_3 & heap_bh30_w77_2 & heap_bh30_w77_1 & heap_bh30_w77_0;
   CompressorIn_bh30_121_213(0) <= heap_bh30_w78_2;
      Compressor_bh30_121: Compressor_14_3
      port map ( R => CompressorOut_bh30_121_121,
                 X0 => CompressorIn_bh30_121_212,
                 X1 => CompressorIn_bh30_121_213);
   heap_bh30_w77_5 <= CompressorOut_bh30_121_121(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w78_3 <= CompressorOut_bh30_121_121(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w79_3 <= CompressorOut_bh30_121_121(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_122_214 <= heap_bh30_w36_11 & heap_bh30_w36_7 & heap_bh30_w36_6 & heap_bh30_w36_5 & heap_bh30_w36_4;
      Compressor_bh30_122: Compressor_5_3
      port map ( R => CompressorOut_bh30_122_122,
                 X0 => CompressorIn_bh30_122_214);
   heap_bh30_w36_13 <= CompressorOut_bh30_122_122(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w37_14 <= CompressorOut_bh30_122_122(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w38_15 <= CompressorOut_bh30_122_122(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_123_215 <= heap_bh30_w22_9 & heap_bh30_w22_5 & heap_bh30_w22_4 & heap_bh30_w22_3;
      Compressor_bh30_123: Compressor_4_3
      port map ( R => CompressorOut_bh30_123_123,
                 X0 => CompressorIn_bh30_123_215);
   heap_bh30_w22_11 <= CompressorOut_bh30_123_123(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w23_13 <= CompressorOut_bh30_123_123(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w24_14 <= CompressorOut_bh30_123_123(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_124_216 <= heap_bh30_w25_6 & heap_bh30_w25_5 & heap_bh30_w25_4 & heap_bh30_w25_3;
      Compressor_bh30_124: Compressor_4_3
      port map ( R => CompressorOut_bh30_124_124,
                 X0 => CompressorIn_bh30_124_216);
   heap_bh30_w25_13 <= CompressorOut_bh30_124_124(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w26_14 <= CompressorOut_bh30_124_124(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w27_14 <= CompressorOut_bh30_124_124(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_125_217 <= heap_bh30_w28_6 & heap_bh30_w28_5 & heap_bh30_w28_4 & heap_bh30_w28_3;
      Compressor_bh30_125: Compressor_4_3
      port map ( R => CompressorOut_bh30_125_125,
                 X0 => CompressorIn_bh30_125_217);
   heap_bh30_w28_13 <= CompressorOut_bh30_125_125(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w29_14 <= CompressorOut_bh30_125_125(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w30_14 <= CompressorOut_bh30_125_125(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_126_218 <= heap_bh30_w31_6 & heap_bh30_w31_5 & heap_bh30_w31_4 & heap_bh30_w31_3;
      Compressor_bh30_126: Compressor_4_3
      port map ( R => CompressorOut_bh30_126_126,
                 X0 => CompressorIn_bh30_126_218);
   heap_bh30_w31_13 <= CompressorOut_bh30_126_126(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w32_14 <= CompressorOut_bh30_126_126(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w33_14 <= CompressorOut_bh30_126_126(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_127_219 <= heap_bh30_w34_6 & heap_bh30_w34_5 & heap_bh30_w34_4 & heap_bh30_w34_3;
      Compressor_bh30_127: Compressor_4_3
      port map ( R => CompressorOut_bh30_127_127,
                 X0 => CompressorIn_bh30_127_219);
   heap_bh30_w34_13 <= CompressorOut_bh30_127_127(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w35_14 <= CompressorOut_bh30_127_127(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w36_14 <= CompressorOut_bh30_127_127(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_128_220 <= heap_bh30_w3_0 & heap_bh30_w3_4 & heap_bh30_w3_3;
   CompressorIn_bh30_128_221 <= heap_bh30_w4_5 & heap_bh30_w4_4;
      Compressor_bh30_128: Compressor_23_3
      port map ( R => CompressorOut_bh30_128_128,
                 X0 => CompressorIn_bh30_128_220,
                 X1 => CompressorIn_bh30_128_221);
   heap_bh30_w3_5 <= CompressorOut_bh30_128_128(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w4_6 <= CompressorOut_bh30_128_128(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w5_7 <= CompressorOut_bh30_128_128(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_129_222 <= heap_bh30_w8_8 & heap_bh30_w8_5 & heap_bh30_w8_4;
   CompressorIn_bh30_129_223 <= heap_bh30_w9_9 & heap_bh30_w9_5;
      Compressor_bh30_129: Compressor_23_3
      port map ( R => CompressorOut_bh30_129_129,
                 X0 => CompressorIn_bh30_129_222,
                 X1 => CompressorIn_bh30_129_223);
   heap_bh30_w8_10 <= CompressorOut_bh30_129_129(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w9_10 <= CompressorOut_bh30_129_129(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w10_9 <= CompressorOut_bh30_129_129(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_130_224 <= heap_bh30_w79_2 & heap_bh30_w79_1 & heap_bh30_w79_0;
   CompressorIn_bh30_130_225 <= heap_bh30_w80_2 & heap_bh30_w80_1;
      Compressor_bh30_130: Compressor_23_3
      port map ( R => CompressorOut_bh30_130_130,
                 X0 => CompressorIn_bh30_130_224,
                 X1 => CompressorIn_bh30_130_225);
   heap_bh30_w79_4 <= CompressorOut_bh30_130_130(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w80_3 <= CompressorOut_bh30_130_130(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w81_3 <= CompressorOut_bh30_130_130(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_131_226 <= heap_bh30_w81_2 & heap_bh30_w81_1 & heap_bh30_w81_0;
   CompressorIn_bh30_131_227 <= heap_bh30_w82_2 & heap_bh30_w82_1;
      Compressor_bh30_131: Compressor_23_3
      port map ( R => CompressorOut_bh30_131_131,
                 X0 => CompressorIn_bh30_131_226,
                 X1 => CompressorIn_bh30_131_227);
   heap_bh30_w81_4 <= CompressorOut_bh30_131_131(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w82_3 <= CompressorOut_bh30_131_131(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w83_3 <= CompressorOut_bh30_131_131(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_132_228 <= heap_bh30_w83_2 & heap_bh30_w83_1 & heap_bh30_w83_0;
   CompressorIn_bh30_132_229 <= heap_bh30_w84_2 & heap_bh30_w84_1;
      Compressor_bh30_132: Compressor_23_3
      port map ( R => CompressorOut_bh30_132_132,
                 X0 => CompressorIn_bh30_132_228,
                 X1 => CompressorIn_bh30_132_229);
   heap_bh30_w83_4 <= CompressorOut_bh30_132_132(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w84_3 <= CompressorOut_bh30_132_132(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w85_3 <= CompressorOut_bh30_132_132(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_133_230 <= heap_bh30_w85_2 & heap_bh30_w85_1 & heap_bh30_w85_0;
   CompressorIn_bh30_133_231 <= heap_bh30_w86_2 & heap_bh30_w86_1;
      Compressor_bh30_133: Compressor_23_3
      port map ( R => CompressorOut_bh30_133_133,
                 X0 => CompressorIn_bh30_133_230,
                 X1 => CompressorIn_bh30_133_231);
   heap_bh30_w85_4 <= CompressorOut_bh30_133_133(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w86_3 <= CompressorOut_bh30_133_133(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w87_3 <= CompressorOut_bh30_133_133(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_134_232 <= heap_bh30_w87_2 & heap_bh30_w87_1 & heap_bh30_w87_0;
   CompressorIn_bh30_134_233 <= heap_bh30_w88_1 & heap_bh30_w88_0;
      Compressor_bh30_134: Compressor_23_3
      port map ( R => CompressorOut_bh30_134_134,
                 X0 => CompressorIn_bh30_134_232,
                 X1 => CompressorIn_bh30_134_233);
   heap_bh30_w87_4 <= CompressorOut_bh30_134_134(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w88_2 <= CompressorOut_bh30_134_134(1); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w89_2 <= CompressorOut_bh30_134_134(2); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_135_234 <= heap_bh30_w5_6 & heap_bh30_w5_5 & heap_bh30_w5_4;
      Compressor_bh30_135: Compressor_3_2
      port map ( R => CompressorOut_bh30_135_135,
                 X0 => CompressorIn_bh30_135_234);
   heap_bh30_w5_8 <= CompressorOut_bh30_135_135(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w6_9 <= CompressorOut_bh30_135_135(1); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_136_235 <= heap_bh30_w10_8 & heap_bh30_w10_4 & heap_bh30_w10_3;
      Compressor_bh30_136: Compressor_3_2
      port map ( R => CompressorOut_bh30_136_136,
                 X0 => CompressorIn_bh30_136_235);
   heap_bh30_w10_10 <= CompressorOut_bh30_136_136(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w11_11 <= CompressorOut_bh30_136_136(1); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_137_236 <= heap_bh30_w15_6 & heap_bh30_w15_5 & heap_bh30_w15_4;
      Compressor_bh30_137: Compressor_3_2
      port map ( R => CompressorOut_bh30_137_137,
                 X0 => CompressorIn_bh30_137_236);
   heap_bh30_w15_13 <= CompressorOut_bh30_137_137(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w16_12 <= CompressorOut_bh30_137_137(1); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_138_237 <= heap_bh30_w18_6 & heap_bh30_w18_5 & heap_bh30_w18_4;
      Compressor_bh30_138: Compressor_3_2
      port map ( R => CompressorOut_bh30_138_138,
                 X0 => CompressorIn_bh30_138_237);
   heap_bh30_w18_13 <= CompressorOut_bh30_138_138(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w19_12 <= CompressorOut_bh30_138_138(1); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_139_238 <= heap_bh30_w21_6 & heap_bh30_w21_5 & heap_bh30_w21_4;
      Compressor_bh30_139: Compressor_3_2
      port map ( R => CompressorOut_bh30_139_139,
                 X0 => CompressorIn_bh30_139_238);
   heap_bh30_w21_13 <= CompressorOut_bh30_139_139(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w22_12 <= CompressorOut_bh30_139_139(1); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_140_239 <= heap_bh30_w64_2 & heap_bh30_w64_1 & heap_bh30_w64_0;
      Compressor_bh30_140: Compressor_3_2
      port map ( R => CompressorOut_bh30_140_140,
                 X0 => CompressorIn_bh30_140_239);
   heap_bh30_w64_6 <= CompressorOut_bh30_140_140(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w65_6 <= CompressorOut_bh30_140_140(1); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_141_240 <= heap_bh30_w66_2 & heap_bh30_w66_1 & heap_bh30_w66_0;
      Compressor_bh30_141: Compressor_3_2
      port map ( R => CompressorOut_bh30_141_141,
                 X0 => CompressorIn_bh30_141_240);
   heap_bh30_w66_5 <= CompressorOut_bh30_141_141(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w67_6 <= CompressorOut_bh30_141_141(1); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_142_241 <= heap_bh30_w68_2 & heap_bh30_w68_1 & heap_bh30_w68_0;
      Compressor_bh30_142: Compressor_3_2
      port map ( R => CompressorOut_bh30_142_142,
                 X0 => CompressorIn_bh30_142_241);
   heap_bh30_w68_5 <= CompressorOut_bh30_142_142(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w69_6 <= CompressorOut_bh30_142_142(1); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_143_242 <= heap_bh30_w70_2 & heap_bh30_w70_1 & heap_bh30_w70_0;
      Compressor_bh30_143: Compressor_3_2
      port map ( R => CompressorOut_bh30_143_143,
                 X0 => CompressorIn_bh30_143_242);
   heap_bh30_w70_5 <= CompressorOut_bh30_143_143(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w71_6 <= CompressorOut_bh30_143_143(1); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_144_243 <= heap_bh30_w72_2 & heap_bh30_w72_1 & heap_bh30_w72_0;
      Compressor_bh30_144: Compressor_3_2
      port map ( R => CompressorOut_bh30_144_144,
                 X0 => CompressorIn_bh30_144_243);
   heap_bh30_w72_5 <= CompressorOut_bh30_144_144(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w73_6 <= CompressorOut_bh30_144_144(1); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_145_244 <= heap_bh30_w74_2 & heap_bh30_w74_1 & heap_bh30_w74_0;
      Compressor_bh30_145: Compressor_3_2
      port map ( R => CompressorOut_bh30_145_145,
                 X0 => CompressorIn_bh30_145_244);
   heap_bh30_w74_5 <= CompressorOut_bh30_145_145(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w75_6 <= CompressorOut_bh30_145_145(1); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_146_245 <= heap_bh30_w76_2 & heap_bh30_w76_1 & heap_bh30_w76_0;
      Compressor_bh30_146: Compressor_3_2
      port map ( R => CompressorOut_bh30_146_146,
                 X0 => CompressorIn_bh30_146_245);
   heap_bh30_w76_5 <= CompressorOut_bh30_146_146(0); -- cycle= 0 cp= 2.91772e-09
   heap_bh30_w77_6 <= CompressorOut_bh30_146_146(1); -- cycle= 0 cp= 2.91772e-09

   CompressorIn_bh30_147_246 <= heap_bh30_w24_4 & heap_bh30_w24_14 & heap_bh30_w24_13 & heap_bh30_w24_12;
   CompressorIn_bh30_147_247(0) <= heap_bh30_w25_13;
      Compressor_bh30_147: Compressor_14_3
      port map ( R => CompressorOut_bh30_147_147,
                 X0 => CompressorIn_bh30_147_246,
                 X1 => CompressorIn_bh30_147_247);
   heap_bh30_w24_15 <= CompressorOut_bh30_147_147(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w25_14 <= CompressorOut_bh30_147_147(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w26_15 <= CompressorOut_bh30_147_147(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_148_248 <= heap_bh30_w27_4 & heap_bh30_w27_14 & heap_bh30_w27_13 & heap_bh30_w27_12;
   CompressorIn_bh30_148_249(0) <= heap_bh30_w28_13;
      Compressor_bh30_148: Compressor_14_3
      port map ( R => CompressorOut_bh30_148_148,
                 X0 => CompressorIn_bh30_148_248,
                 X1 => CompressorIn_bh30_148_249);
   heap_bh30_w27_15 <= CompressorOut_bh30_148_148(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w28_14 <= CompressorOut_bh30_148_148(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w29_15 <= CompressorOut_bh30_148_148(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_149_250 <= heap_bh30_w30_4 & heap_bh30_w30_14 & heap_bh30_w30_13 & heap_bh30_w30_12;
   CompressorIn_bh30_149_251(0) <= heap_bh30_w31_13;
      Compressor_bh30_149: Compressor_14_3
      port map ( R => CompressorOut_bh30_149_149,
                 X0 => CompressorIn_bh30_149_250,
                 X1 => CompressorIn_bh30_149_251);
   heap_bh30_w30_15 <= CompressorOut_bh30_149_149(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w31_14 <= CompressorOut_bh30_149_149(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w32_15 <= CompressorOut_bh30_149_149(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_150_252 <= heap_bh30_w33_4 & heap_bh30_w33_14 & heap_bh30_w33_13 & heap_bh30_w33_12;
   CompressorIn_bh30_150_253(0) <= heap_bh30_w34_13;
      Compressor_bh30_150: Compressor_14_3
      port map ( R => CompressorOut_bh30_150_150,
                 X0 => CompressorIn_bh30_150_252,
                 X1 => CompressorIn_bh30_150_253);
   heap_bh30_w33_15 <= CompressorOut_bh30_150_150(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w34_14 <= CompressorOut_bh30_150_150(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w35_15 <= CompressorOut_bh30_150_150(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_151_254 <= heap_bh30_w38_4 & heap_bh30_w38_15 & heap_bh30_w38_14 & heap_bh30_w38_13;
   CompressorIn_bh30_151_255(0) <= heap_bh30_w39_15;
      Compressor_bh30_151: Compressor_14_3
      port map ( R => CompressorOut_bh30_151_151,
                 X0 => CompressorIn_bh30_151_254,
                 X1 => CompressorIn_bh30_151_255);
   heap_bh30_w38_16 <= CompressorOut_bh30_151_151(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w39_16 <= CompressorOut_bh30_151_151(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w40_15 <= CompressorOut_bh30_151_151(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_152_256 <= heap_bh30_w41_4 & heap_bh30_w41_15 & heap_bh30_w41_14 & heap_bh30_w41_13;
   CompressorIn_bh30_152_257(0) <= heap_bh30_w42_15;
      Compressor_bh30_152: Compressor_14_3
      port map ( R => CompressorOut_bh30_152_152,
                 X0 => CompressorIn_bh30_152_256,
                 X1 => CompressorIn_bh30_152_257);
   heap_bh30_w41_16 <= CompressorOut_bh30_152_152(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w42_16 <= CompressorOut_bh30_152_152(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w43_15 <= CompressorOut_bh30_152_152(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_153_258 <= heap_bh30_w44_4 & heap_bh30_w44_15 & heap_bh30_w44_14 & heap_bh30_w44_13;
   CompressorIn_bh30_153_259(0) <= heap_bh30_w45_15;
      Compressor_bh30_153: Compressor_14_3
      port map ( R => CompressorOut_bh30_153_153,
                 X0 => CompressorIn_bh30_153_258,
                 X1 => CompressorIn_bh30_153_259);
   heap_bh30_w44_16 <= CompressorOut_bh30_153_153(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w45_16 <= CompressorOut_bh30_153_153(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w46_15 <= CompressorOut_bh30_153_153(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_154_260 <= heap_bh30_w47_4 & heap_bh30_w47_15 & heap_bh30_w47_14 & heap_bh30_w47_13;
   CompressorIn_bh30_154_261(0) <= heap_bh30_w48_15;
      Compressor_bh30_154: Compressor_14_3
      port map ( R => CompressorOut_bh30_154_154,
                 X0 => CompressorIn_bh30_154_260,
                 X1 => CompressorIn_bh30_154_261);
   heap_bh30_w47_16 <= CompressorOut_bh30_154_154(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w48_16 <= CompressorOut_bh30_154_154(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w49_15 <= CompressorOut_bh30_154_154(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_155_262 <= heap_bh30_w50_4 & heap_bh30_w50_15 & heap_bh30_w50_14 & heap_bh30_w50_13;
   CompressorIn_bh30_155_263(0) <= heap_bh30_w51_15;
      Compressor_bh30_155: Compressor_14_3
      port map ( R => CompressorOut_bh30_155_155,
                 X0 => CompressorIn_bh30_155_262,
                 X1 => CompressorIn_bh30_155_263);
   heap_bh30_w50_16 <= CompressorOut_bh30_155_155(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w51_16 <= CompressorOut_bh30_155_155(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w52_15 <= CompressorOut_bh30_155_155(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_156_264 <= heap_bh30_w53_4 & heap_bh30_w53_15 & heap_bh30_w53_14 & heap_bh30_w53_13;
   CompressorIn_bh30_156_265(0) <= heap_bh30_w54_15;
      Compressor_bh30_156: Compressor_14_3
      port map ( R => CompressorOut_bh30_156_156,
                 X0 => CompressorIn_bh30_156_264,
                 X1 => CompressorIn_bh30_156_265);
   heap_bh30_w53_16 <= CompressorOut_bh30_156_156(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w54_16 <= CompressorOut_bh30_156_156(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w55_15 <= CompressorOut_bh30_156_156(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_157_266 <= heap_bh30_w56_3 & heap_bh30_w56_14 & heap_bh30_w56_13 & heap_bh30_w56_12;
   CompressorIn_bh30_157_267(0) <= heap_bh30_w57_13;
      Compressor_bh30_157: Compressor_14_3
      port map ( R => CompressorOut_bh30_157_157,
                 X0 => CompressorIn_bh30_157_266,
                 X1 => CompressorIn_bh30_157_267);
   heap_bh30_w56_15 <= CompressorOut_bh30_157_157(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w57_14 <= CompressorOut_bh30_157_157(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w58_11 <= CompressorOut_bh30_157_157(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_158_268 <= heap_bh30_w59_1 & heap_bh30_w59_9 & heap_bh30_w59_8 & heap_bh30_w59_7;
   CompressorIn_bh30_158_269(0) <= heap_bh30_w60_8;
      Compressor_bh30_158: Compressor_14_3
      port map ( R => CompressorOut_bh30_158_158,
                 X0 => CompressorIn_bh30_158_268,
                 X1 => CompressorIn_bh30_158_269);
   heap_bh30_w59_10 <= CompressorOut_bh30_158_158(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w60_9 <= CompressorOut_bh30_158_158(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w61_8 <= CompressorOut_bh30_158_158(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_159_270 <= heap_bh30_w61_0 & heap_bh30_w61_7 & heap_bh30_w61_6 & heap_bh30_w61_5;
   CompressorIn_bh30_159_271(0) <= heap_bh30_w62_7;
      Compressor_bh30_159: Compressor_14_3
      port map ( R => CompressorOut_bh30_159_159,
                 X0 => CompressorIn_bh30_159_270,
                 X1 => CompressorIn_bh30_159_271);
   heap_bh30_w61_9 <= CompressorOut_bh30_159_159(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w62_8 <= CompressorOut_bh30_159_159(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w63_8 <= CompressorOut_bh30_159_159(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_160_272 <= heap_bh30_w7_4 & heap_bh30_w7_3 & heap_bh30_w7_8;
   CompressorIn_bh30_160_273 <= heap_bh30_w8_10 & heap_bh30_w8_9;
      Compressor_bh30_160: Compressor_23_3
      port map ( R => CompressorOut_bh30_160_160,
                 X0 => CompressorIn_bh30_160_272,
                 X1 => CompressorIn_bh30_160_273);
   heap_bh30_w7_9 <= CompressorOut_bh30_160_160(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w8_11 <= CompressorOut_bh30_160_160(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w9_11 <= CompressorOut_bh30_160_160(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_161_274 <= heap_bh30_w12_5 & heap_bh30_w12_4 & heap_bh30_w12_10;
   CompressorIn_bh30_161_275 <= heap_bh30_w13_11 & heap_bh30_w13_10;
      Compressor_bh30_161: Compressor_23_3
      port map ( R => CompressorOut_bh30_161_161,
                 X0 => CompressorIn_bh30_161_274,
                 X1 => CompressorIn_bh30_161_275);
   heap_bh30_w12_11 <= CompressorOut_bh30_161_161(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w13_12 <= CompressorOut_bh30_161_161(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w14_13 <= CompressorOut_bh30_161_161(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_162_276 <= heap_bh30_w15_13 & heap_bh30_w15_12 & heap_bh30_w15_11;
   CompressorIn_bh30_162_277 <= heap_bh30_w16_12 & heap_bh30_w16_11;
      Compressor_bh30_162: Compressor_23_3
      port map ( R => CompressorOut_bh30_162_162,
                 X0 => CompressorIn_bh30_162_276,
                 X1 => CompressorIn_bh30_162_277);
   heap_bh30_w15_14 <= CompressorOut_bh30_162_162(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w16_13 <= CompressorOut_bh30_162_162(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w17_13 <= CompressorOut_bh30_162_162(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_163_278 <= heap_bh30_w18_13 & heap_bh30_w18_12 & heap_bh30_w18_11;
   CompressorIn_bh30_163_279 <= heap_bh30_w19_12 & heap_bh30_w19_11;
      Compressor_bh30_163: Compressor_23_3
      port map ( R => CompressorOut_bh30_163_163,
                 X0 => CompressorIn_bh30_163_278,
                 X1 => CompressorIn_bh30_163_279);
   heap_bh30_w18_14 <= CompressorOut_bh30_163_163(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w19_13 <= CompressorOut_bh30_163_163(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w20_13 <= CompressorOut_bh30_163_163(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_164_280 <= heap_bh30_w21_13 & heap_bh30_w21_12 & heap_bh30_w21_11;
   CompressorIn_bh30_164_281 <= heap_bh30_w22_12 & heap_bh30_w22_11;
      Compressor_bh30_164: Compressor_23_3
      port map ( R => CompressorOut_bh30_164_164,
                 X0 => CompressorIn_bh30_164_280,
                 X1 => CompressorIn_bh30_164_281);
   heap_bh30_w21_14 <= CompressorOut_bh30_164_164(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w22_13 <= CompressorOut_bh30_164_164(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w23_14 <= CompressorOut_bh30_164_164(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_165_282 <= heap_bh30_w35_14 & heap_bh30_w35_13 & heap_bh30_w35_12;
   CompressorIn_bh30_165_283 <= heap_bh30_w36_14 & heap_bh30_w36_13;
      Compressor_bh30_165: Compressor_23_3
      port map ( R => CompressorOut_bh30_165_165,
                 X0 => CompressorIn_bh30_165_282,
                 X1 => CompressorIn_bh30_165_283);
   heap_bh30_w35_16 <= CompressorOut_bh30_165_165(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w36_15 <= CompressorOut_bh30_165_165(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w37_15 <= CompressorOut_bh30_165_165(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_166_284 <= heap_bh30_w63_7 & heap_bh30_w63_6 & heap_bh30_w63_5;
   CompressorIn_bh30_166_285 <= heap_bh30_w64_6 & heap_bh30_w64_5;
      Compressor_bh30_166: Compressor_23_3
      port map ( R => CompressorOut_bh30_166_166,
                 X0 => CompressorIn_bh30_166_284,
                 X1 => CompressorIn_bh30_166_285);
   heap_bh30_w63_9 <= CompressorOut_bh30_166_166(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w64_7 <= CompressorOut_bh30_166_166(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w65_7 <= CompressorOut_bh30_166_166(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_167_286 <= heap_bh30_w65_6 & heap_bh30_w65_5 & heap_bh30_w65_4;
   CompressorIn_bh30_167_287 <= heap_bh30_w66_5 & heap_bh30_w66_4;
      Compressor_bh30_167: Compressor_23_3
      port map ( R => CompressorOut_bh30_167_167,
                 X0 => CompressorIn_bh30_167_286,
                 X1 => CompressorIn_bh30_167_287);
   heap_bh30_w65_8 <= CompressorOut_bh30_167_167(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w66_6 <= CompressorOut_bh30_167_167(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w67_7 <= CompressorOut_bh30_167_167(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_168_288 <= heap_bh30_w67_6 & heap_bh30_w67_5 & heap_bh30_w67_4;
   CompressorIn_bh30_168_289 <= heap_bh30_w68_5 & heap_bh30_w68_4;
      Compressor_bh30_168: Compressor_23_3
      port map ( R => CompressorOut_bh30_168_168,
                 X0 => CompressorIn_bh30_168_288,
                 X1 => CompressorIn_bh30_168_289);
   heap_bh30_w67_8 <= CompressorOut_bh30_168_168(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w68_6 <= CompressorOut_bh30_168_168(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w69_7 <= CompressorOut_bh30_168_168(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_169_290 <= heap_bh30_w69_6 & heap_bh30_w69_5 & heap_bh30_w69_4;
   CompressorIn_bh30_169_291 <= heap_bh30_w70_5 & heap_bh30_w70_4;
      Compressor_bh30_169: Compressor_23_3
      port map ( R => CompressorOut_bh30_169_169,
                 X0 => CompressorIn_bh30_169_290,
                 X1 => CompressorIn_bh30_169_291);
   heap_bh30_w69_8 <= CompressorOut_bh30_169_169(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w70_6 <= CompressorOut_bh30_169_169(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w71_7 <= CompressorOut_bh30_169_169(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_170_292 <= heap_bh30_w71_6 & heap_bh30_w71_5 & heap_bh30_w71_4;
   CompressorIn_bh30_170_293 <= heap_bh30_w72_5 & heap_bh30_w72_4;
      Compressor_bh30_170: Compressor_23_3
      port map ( R => CompressorOut_bh30_170_170,
                 X0 => CompressorIn_bh30_170_292,
                 X1 => CompressorIn_bh30_170_293);
   heap_bh30_w71_8 <= CompressorOut_bh30_170_170(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w72_6 <= CompressorOut_bh30_170_170(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w73_7 <= CompressorOut_bh30_170_170(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_171_294 <= heap_bh30_w73_6 & heap_bh30_w73_5 & heap_bh30_w73_4;
   CompressorIn_bh30_171_295 <= heap_bh30_w74_5 & heap_bh30_w74_4;
      Compressor_bh30_171: Compressor_23_3
      port map ( R => CompressorOut_bh30_171_171,
                 X0 => CompressorIn_bh30_171_294,
                 X1 => CompressorIn_bh30_171_295);
   heap_bh30_w73_8 <= CompressorOut_bh30_171_171(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w74_6 <= CompressorOut_bh30_171_171(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w75_7 <= CompressorOut_bh30_171_171(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_172_296 <= heap_bh30_w75_6 & heap_bh30_w75_5 & heap_bh30_w75_4;
   CompressorIn_bh30_172_297 <= heap_bh30_w76_5 & heap_bh30_w76_4;
      Compressor_bh30_172: Compressor_23_3
      port map ( R => CompressorOut_bh30_172_172,
                 X0 => CompressorIn_bh30_172_296,
                 X1 => CompressorIn_bh30_172_297);
   heap_bh30_w75_8 <= CompressorOut_bh30_172_172(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w76_6 <= CompressorOut_bh30_172_172(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w77_7 <= CompressorOut_bh30_172_172(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_173_298 <= heap_bh30_w77_6 & heap_bh30_w77_5 & heap_bh30_w77_4;
   CompressorIn_bh30_173_299 <= heap_bh30_w78_1 & heap_bh30_w78_0;
      Compressor_bh30_173: Compressor_23_3
      port map ( R => CompressorOut_bh30_173_173,
                 X0 => CompressorIn_bh30_173_298,
                 X1 => CompressorIn_bh30_173_299);
   heap_bh30_w77_8 <= CompressorOut_bh30_173_173(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w78_4 <= CompressorOut_bh30_173_173(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w79_5 <= CompressorOut_bh30_173_173(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_174_300 <= heap_bh30_w89_1 & heap_bh30_w89_0 & heap_bh30_w89_2;
   CompressorIn_bh30_174_301 <= heap_bh30_w90_1 & heap_bh30_w90_0;
      Compressor_bh30_174: Compressor_23_3
      port map ( R => CompressorOut_bh30_174_174,
                 X0 => CompressorIn_bh30_174_300,
                 X1 => CompressorIn_bh30_174_301);
   heap_bh30_w89_3 <= CompressorOut_bh30_174_174(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w90_2 <= CompressorOut_bh30_174_174(1); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w91_2 <= CompressorOut_bh30_174_174(2); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_175_302 <= heap_bh30_w26_14 & heap_bh30_w26_13 & heap_bh30_w26_12;
      Compressor_bh30_175: Compressor_3_2
      port map ( R => CompressorOut_bh30_175_175,
                 X0 => CompressorIn_bh30_175_302);
   heap_bh30_w26_16 <= CompressorOut_bh30_175_175(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w27_16 <= CompressorOut_bh30_175_175(1); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_176_303 <= heap_bh30_w29_14 & heap_bh30_w29_13 & heap_bh30_w29_12;
      Compressor_bh30_176: Compressor_3_2
      port map ( R => CompressorOut_bh30_176_176,
                 X0 => CompressorIn_bh30_176_303);
   heap_bh30_w29_16 <= CompressorOut_bh30_176_176(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w30_16 <= CompressorOut_bh30_176_176(1); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_177_304 <= heap_bh30_w32_14 & heap_bh30_w32_13 & heap_bh30_w32_12;
      Compressor_bh30_177: Compressor_3_2
      port map ( R => CompressorOut_bh30_177_177,
                 X0 => CompressorIn_bh30_177_304);
   heap_bh30_w32_16 <= CompressorOut_bh30_177_177(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w33_16 <= CompressorOut_bh30_177_177(1); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_178_305 <= heap_bh30_w37_14 & heap_bh30_w37_13 & heap_bh30_w37_12;
      Compressor_bh30_178: Compressor_3_2
      port map ( R => CompressorOut_bh30_178_178,
                 X0 => CompressorIn_bh30_178_305);
   heap_bh30_w37_16 <= CompressorOut_bh30_178_178(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w38_17 <= CompressorOut_bh30_178_178(1); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_179_306 <= heap_bh30_w40_14 & heap_bh30_w40_13 & heap_bh30_w40_12;
      Compressor_bh30_179: Compressor_3_2
      port map ( R => CompressorOut_bh30_179_179,
                 X0 => CompressorIn_bh30_179_306);
   heap_bh30_w40_16 <= CompressorOut_bh30_179_179(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w41_17 <= CompressorOut_bh30_179_179(1); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_180_307 <= heap_bh30_w43_14 & heap_bh30_w43_13 & heap_bh30_w43_12;
      Compressor_bh30_180: Compressor_3_2
      port map ( R => CompressorOut_bh30_180_180,
                 X0 => CompressorIn_bh30_180_307);
   heap_bh30_w43_16 <= CompressorOut_bh30_180_180(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w44_17 <= CompressorOut_bh30_180_180(1); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_181_308 <= heap_bh30_w46_14 & heap_bh30_w46_13 & heap_bh30_w46_12;
      Compressor_bh30_181: Compressor_3_2
      port map ( R => CompressorOut_bh30_181_181,
                 X0 => CompressorIn_bh30_181_308);
   heap_bh30_w46_16 <= CompressorOut_bh30_181_181(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w47_17 <= CompressorOut_bh30_181_181(1); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_182_309 <= heap_bh30_w49_14 & heap_bh30_w49_13 & heap_bh30_w49_12;
      Compressor_bh30_182: Compressor_3_2
      port map ( R => CompressorOut_bh30_182_182,
                 X0 => CompressorIn_bh30_182_309);
   heap_bh30_w49_16 <= CompressorOut_bh30_182_182(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w50_17 <= CompressorOut_bh30_182_182(1); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_183_310 <= heap_bh30_w52_14 & heap_bh30_w52_13 & heap_bh30_w52_12;
      Compressor_bh30_183: Compressor_3_2
      port map ( R => CompressorOut_bh30_183_183,
                 X0 => CompressorIn_bh30_183_310);
   heap_bh30_w52_16 <= CompressorOut_bh30_183_183(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w53_17 <= CompressorOut_bh30_183_183(1); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_184_311 <= heap_bh30_w55_14 & heap_bh30_w55_13 & heap_bh30_w55_12;
      Compressor_bh30_184: Compressor_3_2
      port map ( R => CompressorOut_bh30_184_184,
                 X0 => CompressorIn_bh30_184_311);
   heap_bh30_w55_16 <= CompressorOut_bh30_184_184(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w56_16 <= CompressorOut_bh30_184_184(1); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_185_312 <= heap_bh30_w58_10 & heap_bh30_w58_9 & heap_bh30_w58_8;
      Compressor_bh30_185: Compressor_3_2
      port map ( R => CompressorOut_bh30_185_185,
                 X0 => CompressorIn_bh30_185_312);
   heap_bh30_w58_12 <= CompressorOut_bh30_185_185(0); -- cycle= 0 cp= 3.44844e-09
   heap_bh30_w59_11 <= CompressorOut_bh30_185_185(1); -- cycle= 0 cp= 3.44844e-09

   CompressorIn_bh30_186_313 <= heap_bh30_w9_4 & heap_bh30_w9_10 & heap_bh30_w9_11;
   CompressorIn_bh30_186_314 <= heap_bh30_w10_10 & heap_bh30_w10_9;
      Compressor_bh30_186: Compressor_23_3
      port map ( R => CompressorOut_bh30_186_186,
                 X0 => CompressorIn_bh30_186_313,
                 X1 => CompressorIn_bh30_186_314);
   heap_bh30_w9_12 <= CompressorOut_bh30_186_186(0); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w10_11 <= CompressorOut_bh30_186_186(1); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w11_12 <= CompressorOut_bh30_186_186(2); -- cycle= 0 cp= 3.97916e-09

   CompressorIn_bh30_187_315 <= heap_bh30_w25_12 & heap_bh30_w25_11 & heap_bh30_w25_14;
   CompressorIn_bh30_187_316 <= heap_bh30_w26_16 & heap_bh30_w26_15;
      Compressor_bh30_187: Compressor_23_3
      port map ( R => CompressorOut_bh30_187_187,
                 X0 => CompressorIn_bh30_187_315,
                 X1 => CompressorIn_bh30_187_316);
   heap_bh30_w25_15 <= CompressorOut_bh30_187_187(0); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w26_17 <= CompressorOut_bh30_187_187(1); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w27_17 <= CompressorOut_bh30_187_187(2); -- cycle= 0 cp= 3.97916e-09

   CompressorIn_bh30_188_317 <= heap_bh30_w28_12 & heap_bh30_w28_11 & heap_bh30_w28_14;
   CompressorIn_bh30_188_318 <= heap_bh30_w29_16 & heap_bh30_w29_15;
      Compressor_bh30_188: Compressor_23_3
      port map ( R => CompressorOut_bh30_188_188,
                 X0 => CompressorIn_bh30_188_317,
                 X1 => CompressorIn_bh30_188_318);
   heap_bh30_w28_15 <= CompressorOut_bh30_188_188(0); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w29_17 <= CompressorOut_bh30_188_188(1); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w30_17 <= CompressorOut_bh30_188_188(2); -- cycle= 0 cp= 3.97916e-09

   CompressorIn_bh30_189_319 <= heap_bh30_w31_12 & heap_bh30_w31_11 & heap_bh30_w31_14;
   CompressorIn_bh30_189_320 <= heap_bh30_w32_16 & heap_bh30_w32_15;
      Compressor_bh30_189: Compressor_23_3
      port map ( R => CompressorOut_bh30_189_189,
                 X0 => CompressorIn_bh30_189_319,
                 X1 => CompressorIn_bh30_189_320);
   heap_bh30_w31_15 <= CompressorOut_bh30_189_189(0); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w32_17 <= CompressorOut_bh30_189_189(1); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w33_17 <= CompressorOut_bh30_189_189(2); -- cycle= 0 cp= 3.97916e-09

   CompressorIn_bh30_190_321 <= heap_bh30_w34_12 & heap_bh30_w34_11 & heap_bh30_w34_14;
   CompressorIn_bh30_190_322 <= heap_bh30_w35_16 & heap_bh30_w35_15;
      Compressor_bh30_190: Compressor_23_3
      port map ( R => CompressorOut_bh30_190_190,
                 X0 => CompressorIn_bh30_190_321,
                 X1 => CompressorIn_bh30_190_322);
   heap_bh30_w34_15 <= CompressorOut_bh30_190_190(0); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w35_17 <= CompressorOut_bh30_190_190(1); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w36_16 <= CompressorOut_bh30_190_190(2); -- cycle= 0 cp= 3.97916e-09

   CompressorIn_bh30_191_323 <= heap_bh30_w39_14 & heap_bh30_w39_13 & heap_bh30_w39_16;
   CompressorIn_bh30_191_324 <= heap_bh30_w40_16 & heap_bh30_w40_15;
      Compressor_bh30_191: Compressor_23_3
      port map ( R => CompressorOut_bh30_191_191,
                 X0 => CompressorIn_bh30_191_323,
                 X1 => CompressorIn_bh30_191_324);
   heap_bh30_w39_17 <= CompressorOut_bh30_191_191(0); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w40_17 <= CompressorOut_bh30_191_191(1); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w41_18 <= CompressorOut_bh30_191_191(2); -- cycle= 0 cp= 3.97916e-09

   CompressorIn_bh30_192_325 <= heap_bh30_w42_14 & heap_bh30_w42_13 & heap_bh30_w42_16;
   CompressorIn_bh30_192_326 <= heap_bh30_w43_16 & heap_bh30_w43_15;
      Compressor_bh30_192: Compressor_23_3
      port map ( R => CompressorOut_bh30_192_192,
                 X0 => CompressorIn_bh30_192_325,
                 X1 => CompressorIn_bh30_192_326);
   heap_bh30_w42_17 <= CompressorOut_bh30_192_192(0); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w43_17 <= CompressorOut_bh30_192_192(1); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w44_18 <= CompressorOut_bh30_192_192(2); -- cycle= 0 cp= 3.97916e-09

   CompressorIn_bh30_193_327 <= heap_bh30_w45_14 & heap_bh30_w45_13 & heap_bh30_w45_16;
   CompressorIn_bh30_193_328 <= heap_bh30_w46_16 & heap_bh30_w46_15;
      Compressor_bh30_193: Compressor_23_3
      port map ( R => CompressorOut_bh30_193_193,
                 X0 => CompressorIn_bh30_193_327,
                 X1 => CompressorIn_bh30_193_328);
   heap_bh30_w45_17 <= CompressorOut_bh30_193_193(0); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w46_17 <= CompressorOut_bh30_193_193(1); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w47_18 <= CompressorOut_bh30_193_193(2); -- cycle= 0 cp= 3.97916e-09

   CompressorIn_bh30_194_329 <= heap_bh30_w48_14 & heap_bh30_w48_13 & heap_bh30_w48_16;
   CompressorIn_bh30_194_330 <= heap_bh30_w49_16 & heap_bh30_w49_15;
      Compressor_bh30_194: Compressor_23_3
      port map ( R => CompressorOut_bh30_194_194,
                 X0 => CompressorIn_bh30_194_329,
                 X1 => CompressorIn_bh30_194_330);
   heap_bh30_w48_17 <= CompressorOut_bh30_194_194(0); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w49_17 <= CompressorOut_bh30_194_194(1); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w50_18 <= CompressorOut_bh30_194_194(2); -- cycle= 0 cp= 3.97916e-09

   CompressorIn_bh30_195_331 <= heap_bh30_w51_14 & heap_bh30_w51_13 & heap_bh30_w51_16;
   CompressorIn_bh30_195_332 <= heap_bh30_w52_16 & heap_bh30_w52_15;
      Compressor_bh30_195: Compressor_23_3
      port map ( R => CompressorOut_bh30_195_195,
                 X0 => CompressorIn_bh30_195_331,
                 X1 => CompressorIn_bh30_195_332);
   heap_bh30_w51_17 <= CompressorOut_bh30_195_195(0); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w52_17 <= CompressorOut_bh30_195_195(1); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w53_18 <= CompressorOut_bh30_195_195(2); -- cycle= 0 cp= 3.97916e-09

   CompressorIn_bh30_196_333 <= heap_bh30_w54_14 & heap_bh30_w54_13 & heap_bh30_w54_16;
   CompressorIn_bh30_196_334 <= heap_bh30_w55_16 & heap_bh30_w55_15;
      Compressor_bh30_196: Compressor_23_3
      port map ( R => CompressorOut_bh30_196_196,
                 X0 => CompressorIn_bh30_196_333,
                 X1 => CompressorIn_bh30_196_334);
   heap_bh30_w54_17 <= CompressorOut_bh30_196_196(0); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w55_17 <= CompressorOut_bh30_196_196(1); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w56_17 <= CompressorOut_bh30_196_196(2); -- cycle= 0 cp= 3.97916e-09

   CompressorIn_bh30_197_335 <= heap_bh30_w57_12 & heap_bh30_w57_11 & heap_bh30_w57_14;
   CompressorIn_bh30_197_336 <= heap_bh30_w58_12 & heap_bh30_w58_11;
      Compressor_bh30_197: Compressor_23_3
      port map ( R => CompressorOut_bh30_197_197,
                 X0 => CompressorIn_bh30_197_335,
                 X1 => CompressorIn_bh30_197_336);
   heap_bh30_w57_15 <= CompressorOut_bh30_197_197(0); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w58_13 <= CompressorOut_bh30_197_197(1); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w59_12 <= CompressorOut_bh30_197_197(2); -- cycle= 0 cp= 3.97916e-09

   CompressorIn_bh30_198_337 <= heap_bh30_w60_7 & heap_bh30_w60_6 & heap_bh30_w60_9;
   CompressorIn_bh30_198_338 <= heap_bh30_w61_9 & heap_bh30_w61_8;
      Compressor_bh30_198: Compressor_23_3
      port map ( R => CompressorOut_bh30_198_198,
                 X0 => CompressorIn_bh30_198_337,
                 X1 => CompressorIn_bh30_198_338);
   heap_bh30_w60_10 <= CompressorOut_bh30_198_198(0); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w61_10 <= CompressorOut_bh30_198_198(1); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w62_9 <= CompressorOut_bh30_198_198(2); -- cycle= 0 cp= 3.97916e-09

   CompressorIn_bh30_199_339 <= heap_bh30_w62_6 & heap_bh30_w62_5 & heap_bh30_w62_8;
   CompressorIn_bh30_199_340 <= heap_bh30_w63_9 & heap_bh30_w63_8;
      Compressor_bh30_199: Compressor_23_3
      port map ( R => CompressorOut_bh30_199_199,
                 X0 => CompressorIn_bh30_199_339,
                 X1 => CompressorIn_bh30_199_340);
   heap_bh30_w62_10 <= CompressorOut_bh30_199_199(0); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w63_10 <= CompressorOut_bh30_199_199(1); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w64_8 <= CompressorOut_bh30_199_199(2); -- cycle= 0 cp= 3.97916e-09

   CompressorIn_bh30_200_341 <= heap_bh30_w79_4 & heap_bh30_w79_3 & heap_bh30_w79_5;
   CompressorIn_bh30_200_342 <= heap_bh30_w80_0 & heap_bh30_w80_3;
      Compressor_bh30_200: Compressor_23_3
      port map ( R => CompressorOut_bh30_200_200,
                 X0 => CompressorIn_bh30_200_341,
                 X1 => CompressorIn_bh30_200_342);
   heap_bh30_w79_6 <= CompressorOut_bh30_200_200(0); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w80_4 <= CompressorOut_bh30_200_200(1); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w81_5 <= CompressorOut_bh30_200_200(2); -- cycle= 0 cp= 3.97916e-09

   CompressorIn_bh30_201_343 <= heap_bh30_w91_1 & heap_bh30_w91_0 & heap_bh30_w91_2;
   CompressorIn_bh30_201_344 <= heap_bh30_w92_1 & heap_bh30_w92_0;
      Compressor_bh30_201: Compressor_23_3
      port map ( R => CompressorOut_bh30_201_201,
                 X0 => CompressorIn_bh30_201_343,
                 X1 => CompressorIn_bh30_201_344);
   heap_bh30_w91_3 <= CompressorOut_bh30_201_201(0); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w92_2 <= CompressorOut_bh30_201_201(1); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w93_2 <= CompressorOut_bh30_201_201(2); -- cycle= 0 cp= 3.97916e-09

   CompressorIn_bh30_202_345 <= heap_bh30_w14_12 & heap_bh30_w14_11 & heap_bh30_w14_13;
   CompressorIn_bh30_202_346(0) <= heap_bh30_w15_14;
      Compressor_bh30_202: Compressor_13_3
      port map ( R => CompressorOut_bh30_202_202,
                 X0 => CompressorIn_bh30_202_345,
                 X1 => CompressorIn_bh30_202_346);
   heap_bh30_w14_14 <= CompressorOut_bh30_202_202(0); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w15_15 <= CompressorOut_bh30_202_202(1); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w16_14 <= CompressorOut_bh30_202_202(2); -- cycle= 0 cp= 3.97916e-09

   CompressorIn_bh30_203_347 <= heap_bh30_w17_12 & heap_bh30_w17_11 & heap_bh30_w17_13;
   CompressorIn_bh30_203_348(0) <= heap_bh30_w18_14;
      Compressor_bh30_203: Compressor_13_3
      port map ( R => CompressorOut_bh30_203_203,
                 X0 => CompressorIn_bh30_203_347,
                 X1 => CompressorIn_bh30_203_348);
   heap_bh30_w17_14 <= CompressorOut_bh30_203_203(0); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w18_15 <= CompressorOut_bh30_203_203(1); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w19_14 <= CompressorOut_bh30_203_203(2); -- cycle= 0 cp= 3.97916e-09

   CompressorIn_bh30_204_349 <= heap_bh30_w20_12 & heap_bh30_w20_11 & heap_bh30_w20_13;
   CompressorIn_bh30_204_350(0) <= heap_bh30_w21_14;
      Compressor_bh30_204: Compressor_13_3
      port map ( R => CompressorOut_bh30_204_204,
                 X0 => CompressorIn_bh30_204_349,
                 X1 => CompressorIn_bh30_204_350);
   heap_bh30_w20_14 <= CompressorOut_bh30_204_204(0); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w21_15 <= CompressorOut_bh30_204_204(1); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w22_14 <= CompressorOut_bh30_204_204(2); -- cycle= 0 cp= 3.97916e-09

   CompressorIn_bh30_205_351 <= heap_bh30_w23_13 & heap_bh30_w23_12 & heap_bh30_w23_14;
   CompressorIn_bh30_205_352(0) <= heap_bh30_w24_15;
      Compressor_bh30_205: Compressor_13_3
      port map ( R => CompressorOut_bh30_205_205,
                 X0 => CompressorIn_bh30_205_351,
                 X1 => CompressorIn_bh30_205_352);
   heap_bh30_w23_15 <= CompressorOut_bh30_205_205(0); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w24_16 <= CompressorOut_bh30_205_205(1); -- cycle= 0 cp= 3.97916e-09
   heap_bh30_w25_16 <= CompressorOut_bh30_205_205(2); -- cycle= 0 cp= 3.97916e-09

   CompressorIn_bh30_206_353 <= heap_bh30_w36_12 & heap_bh30_w36_15 & heap_bh30_w36_16;
   CompressorIn_bh30_206_354 <= heap_bh30_w37_16 & heap_bh30_w37_15;
      Compressor_bh30_206: Compressor_23_3
      port map ( R => CompressorOut_bh30_206_206,
                 X0 => CompressorIn_bh30_206_353,
                 X1 => CompressorIn_bh30_206_354);
   heap_bh30_w36_17 <= CompressorOut_bh30_206_206(0); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w37_17 <= CompressorOut_bh30_206_206(1); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w38_18 <= CompressorOut_bh30_206_206(2); -- cycle= 0 cp= 4.50988e-09

   CompressorIn_bh30_207_355 <= heap_bh30_w64_4 & heap_bh30_w64_7 & heap_bh30_w64_8;
   CompressorIn_bh30_207_356 <= heap_bh30_w65_8 & heap_bh30_w65_7;
      Compressor_bh30_207: Compressor_23_3
      port map ( R => CompressorOut_bh30_207_207,
                 X0 => CompressorIn_bh30_207_355,
                 X1 => CompressorIn_bh30_207_356);
   heap_bh30_w64_9 <= CompressorOut_bh30_207_207(0); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w65_9 <= CompressorOut_bh30_207_207(1); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w66_7 <= CompressorOut_bh30_207_207(2); -- cycle= 0 cp= 4.50988e-09

   CompressorIn_bh30_208_357 <= heap_bh30_w81_4 & heap_bh30_w81_3 & heap_bh30_w81_5;
   CompressorIn_bh30_208_358 <= heap_bh30_w82_0 & heap_bh30_w82_3;
      Compressor_bh30_208: Compressor_23_3
      port map ( R => CompressorOut_bh30_208_208,
                 X0 => CompressorIn_bh30_208_357,
                 X1 => CompressorIn_bh30_208_358);
   heap_bh30_w81_6 <= CompressorOut_bh30_208_208(0); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w82_4 <= CompressorOut_bh30_208_208(1); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w83_5 <= CompressorOut_bh30_208_208(2); -- cycle= 0 cp= 4.50988e-09

   CompressorIn_bh30_209_359 <= heap_bh30_w93_1 & heap_bh30_w93_0 & heap_bh30_w93_2;
   CompressorIn_bh30_209_360 <= heap_bh30_w94_1 & heap_bh30_w94_0;
      Compressor_bh30_209: Compressor_23_3
      port map ( R => CompressorOut_bh30_209_209,
                 X0 => CompressorIn_bh30_209_359,
                 X1 => CompressorIn_bh30_209_360);
   heap_bh30_w93_3 <= CompressorOut_bh30_209_209(0); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w94_2 <= CompressorOut_bh30_209_209(1); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w95_1 <= CompressorOut_bh30_209_209(2); -- cycle= 0 cp= 4.50988e-09

   CompressorIn_bh30_210_361 <= heap_bh30_w11_11 & heap_bh30_w11_10 & heap_bh30_w11_12;
   CompressorIn_bh30_210_362(0) <= heap_bh30_w12_11;
      Compressor_bh30_210: Compressor_13_3
      port map ( R => CompressorOut_bh30_210_210,
                 X0 => CompressorIn_bh30_210_361,
                 X1 => CompressorIn_bh30_210_362);
   heap_bh30_w11_13 <= CompressorOut_bh30_210_210(0); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w12_12 <= CompressorOut_bh30_210_210(1); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w13_13 <= CompressorOut_bh30_210_210(2); -- cycle= 0 cp= 4.50988e-09

   CompressorIn_bh30_211_363 <= heap_bh30_w16_10 & heap_bh30_w16_13 & heap_bh30_w16_14;
   CompressorIn_bh30_211_364(0) <= heap_bh30_w17_14;
      Compressor_bh30_211: Compressor_13_3
      port map ( R => CompressorOut_bh30_211_211,
                 X0 => CompressorIn_bh30_211_363,
                 X1 => CompressorIn_bh30_211_364);
   heap_bh30_w16_15 <= CompressorOut_bh30_211_211(0); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w17_15 <= CompressorOut_bh30_211_211(1); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w18_16 <= CompressorOut_bh30_211_211(2); -- cycle= 0 cp= 4.50988e-09

   CompressorIn_bh30_212_365 <= heap_bh30_w19_10 & heap_bh30_w19_13 & heap_bh30_w19_14;
   CompressorIn_bh30_212_366(0) <= heap_bh30_w20_14;
      Compressor_bh30_212: Compressor_13_3
      port map ( R => CompressorOut_bh30_212_212,
                 X0 => CompressorIn_bh30_212_365,
                 X1 => CompressorIn_bh30_212_366);
   heap_bh30_w19_15 <= CompressorOut_bh30_212_212(0); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w20_15 <= CompressorOut_bh30_212_212(1); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w21_16 <= CompressorOut_bh30_212_212(2); -- cycle= 0 cp= 4.50988e-09

   CompressorIn_bh30_213_367 <= heap_bh30_w22_10 & heap_bh30_w22_13 & heap_bh30_w22_14;
   CompressorIn_bh30_213_368(0) <= heap_bh30_w23_15;
      Compressor_bh30_213: Compressor_13_3
      port map ( R => CompressorOut_bh30_213_213,
                 X0 => CompressorIn_bh30_213_367,
                 X1 => CompressorIn_bh30_213_368);
   heap_bh30_w22_15 <= CompressorOut_bh30_213_213(0); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w23_16 <= CompressorOut_bh30_213_213(1); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w24_17 <= CompressorOut_bh30_213_213(2); -- cycle= 0 cp= 4.50988e-09

   CompressorIn_bh30_214_369 <= heap_bh30_w27_16 & heap_bh30_w27_15 & heap_bh30_w27_17;
   CompressorIn_bh30_214_370(0) <= heap_bh30_w28_15;
      Compressor_bh30_214: Compressor_13_3
      port map ( R => CompressorOut_bh30_214_214,
                 X0 => CompressorIn_bh30_214_369,
                 X1 => CompressorIn_bh30_214_370);
   heap_bh30_w27_18 <= CompressorOut_bh30_214_214(0); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w28_16 <= CompressorOut_bh30_214_214(1); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w29_18 <= CompressorOut_bh30_214_214(2); -- cycle= 0 cp= 4.50988e-09

   CompressorIn_bh30_215_371 <= heap_bh30_w30_16 & heap_bh30_w30_15 & heap_bh30_w30_17;
   CompressorIn_bh30_215_372(0) <= heap_bh30_w31_15;
      Compressor_bh30_215: Compressor_13_3
      port map ( R => CompressorOut_bh30_215_215,
                 X0 => CompressorIn_bh30_215_371,
                 X1 => CompressorIn_bh30_215_372);
   heap_bh30_w30_18 <= CompressorOut_bh30_215_215(0); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w31_16 <= CompressorOut_bh30_215_215(1); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w32_18 <= CompressorOut_bh30_215_215(2); -- cycle= 0 cp= 4.50988e-09

   CompressorIn_bh30_216_373 <= heap_bh30_w33_16 & heap_bh30_w33_15 & heap_bh30_w33_17;
   CompressorIn_bh30_216_374(0) <= heap_bh30_w34_15;
      Compressor_bh30_216: Compressor_13_3
      port map ( R => CompressorOut_bh30_216_216,
                 X0 => CompressorIn_bh30_216_373,
                 X1 => CompressorIn_bh30_216_374);
   heap_bh30_w33_18 <= CompressorOut_bh30_216_216(0); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w34_16 <= CompressorOut_bh30_216_216(1); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w35_18 <= CompressorOut_bh30_216_216(2); -- cycle= 0 cp= 4.50988e-09

   CompressorIn_bh30_217_375 <= heap_bh30_w41_17 & heap_bh30_w41_16 & heap_bh30_w41_18;
   CompressorIn_bh30_217_376(0) <= heap_bh30_w42_17;
      Compressor_bh30_217: Compressor_13_3
      port map ( R => CompressorOut_bh30_217_217,
                 X0 => CompressorIn_bh30_217_375,
                 X1 => CompressorIn_bh30_217_376);
   heap_bh30_w41_19 <= CompressorOut_bh30_217_217(0); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w42_18 <= CompressorOut_bh30_217_217(1); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w43_18 <= CompressorOut_bh30_217_217(2); -- cycle= 0 cp= 4.50988e-09

   CompressorIn_bh30_218_377 <= heap_bh30_w44_17 & heap_bh30_w44_16 & heap_bh30_w44_18;
   CompressorIn_bh30_218_378(0) <= heap_bh30_w45_17;
      Compressor_bh30_218: Compressor_13_3
      port map ( R => CompressorOut_bh30_218_218,
                 X0 => CompressorIn_bh30_218_377,
                 X1 => CompressorIn_bh30_218_378);
   heap_bh30_w44_19 <= CompressorOut_bh30_218_218(0); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w45_18 <= CompressorOut_bh30_218_218(1); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w46_18 <= CompressorOut_bh30_218_218(2); -- cycle= 0 cp= 4.50988e-09

   CompressorIn_bh30_219_379 <= heap_bh30_w47_17 & heap_bh30_w47_16 & heap_bh30_w47_18;
   CompressorIn_bh30_219_380(0) <= heap_bh30_w48_17;
      Compressor_bh30_219: Compressor_13_3
      port map ( R => CompressorOut_bh30_219_219,
                 X0 => CompressorIn_bh30_219_379,
                 X1 => CompressorIn_bh30_219_380);
   heap_bh30_w47_19 <= CompressorOut_bh30_219_219(0); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w48_18 <= CompressorOut_bh30_219_219(1); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w49_18 <= CompressorOut_bh30_219_219(2); -- cycle= 0 cp= 4.50988e-09

   CompressorIn_bh30_220_381 <= heap_bh30_w50_17 & heap_bh30_w50_16 & heap_bh30_w50_18;
   CompressorIn_bh30_220_382(0) <= heap_bh30_w51_17;
      Compressor_bh30_220: Compressor_13_3
      port map ( R => CompressorOut_bh30_220_220,
                 X0 => CompressorIn_bh30_220_381,
                 X1 => CompressorIn_bh30_220_382);
   heap_bh30_w50_19 <= CompressorOut_bh30_220_220(0); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w51_18 <= CompressorOut_bh30_220_220(1); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w52_18 <= CompressorOut_bh30_220_220(2); -- cycle= 0 cp= 4.50988e-09

   CompressorIn_bh30_221_383 <= heap_bh30_w53_17 & heap_bh30_w53_16 & heap_bh30_w53_18;
   CompressorIn_bh30_221_384(0) <= heap_bh30_w54_17;
      Compressor_bh30_221: Compressor_13_3
      port map ( R => CompressorOut_bh30_221_221,
                 X0 => CompressorIn_bh30_221_383,
                 X1 => CompressorIn_bh30_221_384);
   heap_bh30_w53_19 <= CompressorOut_bh30_221_221(0); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w54_18 <= CompressorOut_bh30_221_221(1); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w55_18 <= CompressorOut_bh30_221_221(2); -- cycle= 0 cp= 4.50988e-09

   CompressorIn_bh30_222_385 <= heap_bh30_w56_16 & heap_bh30_w56_15 & heap_bh30_w56_17;
   CompressorIn_bh30_222_386(0) <= heap_bh30_w57_15;
      Compressor_bh30_222: Compressor_13_3
      port map ( R => CompressorOut_bh30_222_222,
                 X0 => CompressorIn_bh30_222_385,
                 X1 => CompressorIn_bh30_222_386);
   heap_bh30_w56_18 <= CompressorOut_bh30_222_222(0); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w57_16 <= CompressorOut_bh30_222_222(1); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w58_14 <= CompressorOut_bh30_222_222(2); -- cycle= 0 cp= 4.50988e-09

   CompressorIn_bh30_223_387 <= heap_bh30_w59_11 & heap_bh30_w59_10 & heap_bh30_w59_12;
   CompressorIn_bh30_223_388(0) <= heap_bh30_w60_10;
      Compressor_bh30_223: Compressor_13_3
      port map ( R => CompressorOut_bh30_223_223,
                 X0 => CompressorIn_bh30_223_387,
                 X1 => CompressorIn_bh30_223_388);
   heap_bh30_w59_13 <= CompressorOut_bh30_223_223(0); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w60_11 <= CompressorOut_bh30_223_223(1); -- cycle= 0 cp= 4.50988e-09
   heap_bh30_w61_11 <= CompressorOut_bh30_223_223(2); -- cycle= 0 cp= 4.50988e-09

   CompressorIn_bh30_224_389 <= heap_bh30_w83_4 & heap_bh30_w83_3 & heap_bh30_w83_5;
   CompressorIn_bh30_224_390 <= heap_bh30_w84_0 & heap_bh30_w84_3;
      Compressor_bh30_224: Compressor_23_3
      port map ( R => CompressorOut_bh30_224_224,
                 X0 => CompressorIn_bh30_224_389,
                 X1 => CompressorIn_bh30_224_390);
   heap_bh30_w83_6 <= CompressorOut_bh30_224_224(0); -- cycle= 0 cp= 5.0406e-09
   heap_bh30_w84_4 <= CompressorOut_bh30_224_224(1); -- cycle= 0 cp= 5.0406e-09
   heap_bh30_w85_5 <= CompressorOut_bh30_224_224(2); -- cycle= 0 cp= 5.0406e-09

   CompressorIn_bh30_225_391 <= heap_bh30_w38_17 & heap_bh30_w38_16 & heap_bh30_w38_18;
   CompressorIn_bh30_225_392(0) <= heap_bh30_w39_17;
      Compressor_bh30_225: Compressor_13_3
      port map ( R => CompressorOut_bh30_225_225,
                 X0 => CompressorIn_bh30_225_391,
                 X1 => CompressorIn_bh30_225_392);
   heap_bh30_w38_19 <= CompressorOut_bh30_225_225(0); -- cycle= 0 cp= 5.0406e-09
   heap_bh30_w39_18 <= CompressorOut_bh30_225_225(1); -- cycle= 0 cp= 5.0406e-09
   heap_bh30_w40_18 <= CompressorOut_bh30_225_225(2); -- cycle= 0 cp= 5.0406e-09

   CompressorIn_bh30_226_393 <= heap_bh30_w85_4 & heap_bh30_w85_3 & heap_bh30_w85_5;
   CompressorIn_bh30_226_394 <= heap_bh30_w86_0 & heap_bh30_w86_3;
      Compressor_bh30_226: Compressor_23_3
      port map ( R => CompressorOut_bh30_226_226,
                 X0 => CompressorIn_bh30_226_393,
                 X1 => CompressorIn_bh30_226_394);
   heap_bh30_w85_6 <= CompressorOut_bh30_226_226(0); -- cycle= 0 cp= 5.57132e-09
   heap_bh30_w86_4 <= CompressorOut_bh30_226_226(1); -- cycle= 0 cp= 5.57132e-09
   heap_bh30_w87_5 <= CompressorOut_bh30_226_226(2); -- cycle= 0 cp= 5.57132e-09

   CompressorIn_bh30_227_395 <= heap_bh30_w87_4 & heap_bh30_w87_3 & heap_bh30_w87_5;
   CompressorIn_bh30_227_396(0) <= heap_bh30_w88_2;
      Compressor_bh30_227: Compressor_13_3
      port map ( R => CompressorOut_bh30_227_227,
                 X0 => CompressorIn_bh30_227_395,
                 X1 => CompressorIn_bh30_227_396);
   heap_bh30_w87_6 <= CompressorOut_bh30_227_227(0); -- cycle= 0 cp= 6.10204e-09
   heap_bh30_w88_3 <= CompressorOut_bh30_227_227(1); -- cycle= 0 cp= 6.10204e-09
   heap_bh30_w89_4 <= CompressorOut_bh30_227_227(2); -- cycle= 0 cp= 6.10204e-09
   finalAdderIn0_bh30 <= "0" & heap_bh30_w111_0 & heap_bh30_w110_0 & heap_bh30_w109_0 & heap_bh30_w108_0 & heap_bh30_w107_0 & heap_bh30_w106_0 & heap_bh30_w105_0 & heap_bh30_w104_0 & heap_bh30_w103_0 & heap_bh30_w102_0 & heap_bh30_w101_0 & heap_bh30_w100_0 & heap_bh30_w99_0 & heap_bh30_w98_0 & heap_bh30_w97_0 & heap_bh30_w96_0 & heap_bh30_w95_0 & heap_bh30_w94_2 & heap_bh30_w93_3 & heap_bh30_w92_2 & heap_bh30_w91_3 & heap_bh30_w90_2 & heap_bh30_w89_3 & heap_bh30_w88_3 & heap_bh30_w87_6 & heap_bh30_w86_4 & heap_bh30_w85_6 & heap_bh30_w84_4 & heap_bh30_w83_6 & heap_bh30_w82_4 & heap_bh30_w81_6 & heap_bh30_w80_4 & heap_bh30_w79_6 & heap_bh30_w78_3 & heap_bh30_w77_8 & heap_bh30_w76_6 & heap_bh30_w75_8 & heap_bh30_w74_6 & heap_bh30_w73_8 & heap_bh30_w72_6 & heap_bh30_w71_8 & heap_bh30_w70_6 & heap_bh30_w69_8 & heap_bh30_w68_6 & heap_bh30_w67_8 & heap_bh30_w66_6 & heap_bh30_w65_9 & heap_bh30_w64_9 & heap_bh30_w63_10 & heap_bh30_w62_10 & heap_bh30_w61_10 & heap_bh30_w60_11 & heap_bh30_w59_13 & heap_bh30_w58_13 & heap_bh30_w57_16 & heap_bh30_w56_18 & heap_bh30_w55_17 & heap_bh30_w54_18 & heap_bh30_w53_19 & heap_bh30_w52_17 & heap_bh30_w51_18 & heap_bh30_w50_19 & heap_bh30_w49_17 & heap_bh30_w48_18 & heap_bh30_w47_19 & heap_bh30_w46_17 & heap_bh30_w45_18 & heap_bh30_w44_19 & heap_bh30_w43_17 & heap_bh30_w42_18 & heap_bh30_w41_19 & heap_bh30_w40_17 & heap_bh30_w39_18 & heap_bh30_w38_19 & heap_bh30_w37_17 & heap_bh30_w36_17 & heap_bh30_w35_17 & heap_bh30_w34_16 & heap_bh30_w33_18 & heap_bh30_w32_17 & heap_bh30_w31_16 & heap_bh30_w30_18 & heap_bh30_w29_17 & heap_bh30_w28_16 & heap_bh30_w27_18 & heap_bh30_w26_17 & heap_bh30_w25_16 & heap_bh30_w24_16 & heap_bh30_w23_16 & heap_bh30_w22_15 & heap_bh30_w21_15 & heap_bh30_w20_15 & heap_bh30_w19_15 & heap_bh30_w18_15 & heap_bh30_w17_15 & heap_bh30_w16_15 & heap_bh30_w15_15 & heap_bh30_w14_14 & heap_bh30_w13_12 & heap_bh30_w12_12 & heap_bh30_w11_13 & heap_bh30_w10_11 & heap_bh30_w9_12 & heap_bh30_w8_11 & heap_bh30_w7_9 & heap_bh30_w6_9 & heap_bh30_w5_8 & heap_bh30_w4_3 & heap_bh30_w3_5 & heap_bh30_w2_4 & heap_bh30_w1_0 & heap_bh30_w0_0;
   finalAdderIn1_bh30 <= "0" & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & heap_bh30_w95_1 & '0' & '0' & '0' & '0' & '0' & heap_bh30_w89_4 & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & '0' & heap_bh30_w78_4 & heap_bh30_w77_7 & '0' & heap_bh30_w75_7 & '0' & heap_bh30_w73_7 & '0' & heap_bh30_w71_7 & '0' & heap_bh30_w69_7 & '0' & heap_bh30_w67_7 & heap_bh30_w66_7 & '0' & '0' & '0' & heap_bh30_w62_9 & heap_bh30_w61_11 & '0' & '0' & heap_bh30_w58_14 & '0' & '0' & heap_bh30_w55_18 & '0' & '0' & heap_bh30_w52_18 & '0' & '0' & heap_bh30_w49_18 & '0' & '0' & heap_bh30_w46_18 & '0' & '0' & heap_bh30_w43_18 & '0' & '0' & heap_bh30_w40_18 & '0' & '0' & '0' & '0' & heap_bh30_w35_18 & '0' & '0' & heap_bh30_w32_18 & '0' & '0' & heap_bh30_w29_18 & '0' & '0' & '0' & heap_bh30_w25_15 & heap_bh30_w24_17 & '0' & '0' & heap_bh30_w21_16 & '0' & '0' & heap_bh30_w18_16 & '0' & '0' & '0' & '0' & heap_bh30_w13_13 & '0' & '0' & '0' & '0' & '0' & '0' & heap_bh30_w6_8 & heap_bh30_w5_7 & heap_bh30_w4_6 & '0' & heap_bh30_w2_3 & heap_bh30_w1_1 & heap_bh30_w0_1;
   finalAdderCin_bh30 <= '0';
      Adder_final30_0: IntAdder_113_f400_uid580
      port map ( Cin => finalAdderCin_bh30,
                 R => finalAdderOut_bh30,
                 X => finalAdderIn0_bh30,
                 Y => finalAdderIn1_bh30);
   -- concatenate all the compressed chunks
   CompressionResult30 <= finalAdderOut_bh30;
   -- End of code generated by BitHeap::generateCompressorVHDL
   R <= CompressionResult30(111 downto 0);
end architecture;

--------------------------------------------------------------------------------
--                   RightShifter_120_by_max_65_comb_uid590
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Bogdan Pasca, Florent de Dinechin (2008-2011)
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity RightShifter_120_by_max_65_comb_uid590 is
   port ( X : in  std_logic_vector(119 downto 0);
          S : in  std_logic_vector(6 downto 0);
          R : out  std_logic_vector(184 downto 0)   );
end entity;

architecture arch of RightShifter_120_by_max_65_comb_uid590 is
signal level0 :  std_logic_vector(119 downto 0);
signal ps :  std_logic_vector(6 downto 0);
signal level1 :  std_logic_vector(120 downto 0);
signal level2 :  std_logic_vector(122 downto 0);
signal level3 :  std_logic_vector(126 downto 0);
signal level4 :  std_logic_vector(134 downto 0);
signal level5 :  std_logic_vector(150 downto 0);
signal level6 :  std_logic_vector(182 downto 0);
signal level7 :  std_logic_vector(246 downto 0);
begin
   level0<= X;
   ps<= S;
   level1<=  (0 downto 0 => '0') & level0 when ps(0) = '1' else    level0 & (0 downto 0 => '0');
   level2<=  (1 downto 0 => '0') & level1 when ps(1) = '1' else    level1 & (1 downto 0 => '0');
   level3<=  (3 downto 0 => '0') & level2 when ps(2) = '1' else    level2 & (3 downto 0 => '0');
   level4<=  (7 downto 0 => '0') & level3 when ps(3) = '1' else    level3 & (7 downto 0 => '0');
   level5<=  (15 downto 0 => '0') & level4 when ps(4) = '1' else    level4 & (15 downto 0 => '0');
   level6<=  (31 downto 0 => '0') & level5 when ps(5) = '1' else    level5 & (31 downto 0 => '0');
   level7<=  (63 downto 0 => '0') & level6 when ps(6) = '1' else    level6 & (63 downto 0 => '0');
   R <= level7(246 downto 62);
end architecture;

--------------------------------------------------------------------------------
--                          PositMult_65_7_comb_uid2
-- This operator is part of the Infinite Virtual Library FloPoCoLib
-- All rights reserved 
-- Authors: Raul Murillo, 2019
--------------------------------------------------------------------------------
-- combinatorial

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;
library std;
use std.textio.all;
library work;

entity PositMult_65_7_comb_uid2 is
   port ( InputA : in  std_logic_vector(64 downto 0);
          InputB : in  std_logic_vector(64 downto 0);
          Output : out  std_logic_vector(64 downto 0)   );
end entity;

architecture arch of PositMult_65_7_comb_uid2 is
   component PositDecoder_65_7_comb_uid4 is
      port ( Input : in  std_logic_vector(64 downto 0);
             Sign : out  std_logic;
             Reg : out  std_logic_vector(7 downto 0);
             Exp : out  std_logic_vector(6 downto 0);
             Frac : out  std_logic_vector(55 downto 0);
             z : out  std_logic;
             inf : out  std_logic   );
   end component;

   component PositDecoder_65_7_comb_uid16 is
      port ( Input : in  std_logic_vector(64 downto 0);
             Sign : out  std_logic;
             Reg : out  std_logic_vector(7 downto 0);
             Exp : out  std_logic_vector(6 downto 0);
             Frac : out  std_logic_vector(55 downto 0);
             z : out  std_logic;
             inf : out  std_logic   );
   end component;

   component IntMultiplier_UsingDSP_56_56_112_unsigned_comb_uid28 is
      port ( X : in  std_logic_vector(55 downto 0);
             Y : in  std_logic_vector(55 downto 0);
             R : out  std_logic_vector(111 downto 0)   );
   end component;

   component RightShifter_120_by_max_65_comb_uid590 is
      port ( X : in  std_logic_vector(119 downto 0);
             S : in  std_logic_vector(6 downto 0);
             R : out  std_logic_vector(184 downto 0)   );
   end component;

signal sign_A :  std_logic;
signal reg_A :  std_logic_vector(7 downto 0);
signal exp_A :  std_logic_vector(6 downto 0);
signal frac_A :  std_logic_vector(55 downto 0);
signal z_A :  std_logic;
signal inf_A :  std_logic;
signal sign_B :  std_logic;
signal reg_B :  std_logic_vector(7 downto 0);
signal exp_B :  std_logic_vector(6 downto 0);
signal frac_B :  std_logic_vector(55 downto 0);
signal z_B :  std_logic;
signal inf_B :  std_logic;
signal sf_A :  std_logic_vector(14 downto 0);
signal sf_B :  std_logic_vector(14 downto 0);
signal sign :  std_logic;
signal z :  std_logic;
signal inf :  std_logic;
signal frac_mult :  std_logic_vector(111 downto 0);
signal ovf_m :  std_logic;
signal normFrac :  std_logic_vector(112 downto 0);
signal sf_mult :  std_logic_vector(15 downto 0);
signal sf_sign :  std_logic;
signal nzero :  std_logic;
signal ExpBits :  std_logic_vector(6 downto 0);
signal RegimeAns_tmp :  std_logic_vector(6 downto 0);
signal RegimeAns :  std_logic_vector(6 downto 0);
signal ovf_reg :  std_logic;
signal FinalRegime :  std_logic_vector(6 downto 0);
signal ovf_regF :  std_logic;
signal FinalExp :  std_logic_vector(6 downto 0);
signal tmp1 :  std_logic_vector(119 downto 0);
signal tmp2 :  std_logic_vector(119 downto 0);
signal shift_neg :  std_logic_vector(6 downto 0);
signal shift_pos :  std_logic_vector(6 downto 0);
signal shifter_in :  std_logic_vector(119 downto 0);
signal shifter_S :  std_logic_vector(6 downto 0);
signal shifter_out :  std_logic_vector(184 downto 0);
signal tmp_ans :  std_logic_vector(63 downto 0);
signal LSB :  std_logic;
signal G :  std_logic;
signal R :  std_logic;
signal S :  std_logic;
signal round :  std_logic;
begin
------------------------------- Data Extraction -------------------------------
   decoderA: PositDecoder_65_7_comb_uid4
      port map ( Exp => exp_A,
                 Frac => frac_A,
                 Input => InputA,
                 Reg => reg_A,
                 Sign => sign_A,
                 inf => inf_A,
                 z => z_A);
   decoderB: PositDecoder_65_7_comb_uid16
      port map ( Exp => exp_B,
                 Frac => frac_B,
                 Input => InputB,
                 Reg => reg_B,
                 Sign => sign_B,
                 inf => inf_B,
                 z => z_B);
   -- Gather scale factors
   sf_A <= reg_A & exp_A;
   sf_B <= reg_B & exp_B;
---------------------- Sign and Special Cases Computation ----------------------
   sign <= sign_A XOR sign_B;
   z <= z_A OR z_B;
   inf <= inf_A OR inf_B;
--------------- Multiply the fractions, add the exponent values ---------------
   mult: IntMultiplier_UsingDSP_56_56_112_unsigned_comb_uid28
      port map ( R => frac_mult,
                 X => frac_A,
                 Y => frac_B);
   -- Adjust for overflow
   ovf_m <= frac_mult(frac_mult'high);
   normFrac <= frac_mult & '0' when ovf_m = '0' else '0' & frac_mult;
   sf_mult <= (sf_A(sf_A'high) & sf_A) + (sf_B(sf_B'high) & sf_B) + ovf_m;
   sf_sign <= sf_mult(sf_mult'high);
---------------------- Compute Regime and Exponent value ----------------------
   nzero <= '0' when frac_mult = 0 else '1';
   -- Unpack scaling factors
   ExpBits <= sf_mult(6 downto 0);
   RegimeAns_tmp <= sf_mult(13 downto 7);
   -- Get Regime's absolute value
   RegimeAns <= (NOT RegimeAns_tmp)+1 when sf_sign = '1' else RegimeAns_tmp;
   -- Check for Regime overflow
   ovf_reg <= RegimeAns(RegimeAns'high);
   FinalRegime <= '0' & "111111" when ovf_reg = '1' else RegimeAns;
   ovf_regF <= '1' when FinalRegime = ('0' & "111111") else '0';
   FinalExp <= "0000000" when ((ovf_reg = '1') OR (ovf_regF = '1') OR (nzero='0')) else ExpBits;
------------------------------- Packing Stage 1 -------------------------------
   tmp1 <= nzero & '0' & FinalExp & normFrac(110 downto 0);
   tmp2 <= '0' & nzero & FinalExp & normFrac(110 downto 0);
   shift_neg <= FinalRegime - 2 when (ovf_regF = '1') else FinalRegime - 1;
   shift_pos <= FinalRegime - 1 when (ovf_regF = '1') else FinalRegime;
   shifter_in <= tmp2 when sf_sign = '1' else tmp1;
   shifter_S <= shift_neg when sf_sign = '1' else shift_pos;
   RightShifterComponent: RightShifter_120_by_max_65_comb_uid590
      port map ( R => shifter_out,
                 S => shifter_S,
                 X => shifter_in);
   tmp_ans <= shifter_out(184 downto 121);
--------------------- Packing Stage 2 - Unbiased Rounding ---------------------
   LSB <= shifter_out(121);
   G <= shifter_out(120);
   R <= shifter_out(119);
   S <= '0' when shifter_out(118 downto 0) = 0 else '1';
   round <= G AND (LSB OR R OR S) when NOT((ovf_reg OR ovf_regF) = '1') else '0';
   Output <= '1' & "0000000000000000000000000000000000000000000000000000000000000000" when inf = '1' else "00000000000000000000000000000000000000000000000000000000000000000" when z = '1' else '0' & (tmp_ans + round) when sign = '0' else NOT('0' & (tmp_ans + round))+1;
end architecture;

